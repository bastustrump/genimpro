BZh91AY&SYO-R� L_�Ryg����������`+�>$�RP�J��a���ʈ�]w�)�۪֥��jiLMA4�͍)��Q�-�Y�k�sK[lKm����e�&�|}��P��U �dT��� ��0�A� !���ɠ�S�L�H�=i�hb 2a4�i� �EU �12` &��`�����  424   $B4��f)��L$z�S��L���4=C2�@M �i=@ș�S"<MO( �S5v�v�Q���B"(�k).��	�� �n��C� ���uQ�hiǗ�z����N
��{}���#|H������V�;w큛�@���"�� (����@�RJ�t�TuP.R��9�R�A�̪��bi�rأf e�����^�c����a����*��Q�,��;�sEvETI� ���F �}�Lq6`�כ��rqy���9���Fu����<�q���:�,��@$��<���=rDܱY��C�hI4�H�`BU�BuV8��f2���KCAsK�+���t/c5A�e%d�*�b��P�up[�����`��\��-�b���$����<J�i;��ܐ��j�Ef]�Sc0f�t\��!�;�&YޔٮvB�i�-�MڧJ�^��BOK�w/E,����5�.�C�*mP�Y֨$�UXW\ܜ�e�UC2eFK%�H\���P�ANȠ������B���UGg�F	�WZ��]3M��ijPS4�(`�J�<���QVI&rQ����1%\�b*�(.�R#�;�􃒐�".��e+aP�.K�Phu�B��]Hb�,��B����c6�ud&�c�i��*���n-������%j}����wa�ݦi�$K�ؠ�e��ff���|SjD;b�u�m3�ۨ[}H:&;i��R�u+ �(�V�<-u$팱���á' ��K��< ��!`K�v���v1�C��k�oWUb�t���j�t�u��i�HS�'ԞG71�XDɮ8���wn(:�-�N�AB��Kx��In��%�� ����t��|��!q�(Ȏ*K0 �wv[@�cq����ͺډm�mof�A�rkK=x���Zyx몣�8i����q��Qz�Z,���#B���ݱ�bA��}>�)��p�P�#B��%�q^�w�a�AC|���V��� ێS�`��B܌6��?^�����QTm���X�W��za��Ć�U�b_�����v5k��M�+q�v�u�}�eq����� �<0��	�N��X����:ߩc�X�5E�\E� A\�у�ŭ��)�re�F�:�0�-3��}9�n!��D�L�~��m��B�# �
BM~>�.�P&jYY��W�X7�ĞX,B��]�-�.����� U��_�Y�DTR��#�D@t�DCӕ@�`�y��� &A�ʪ\�P��,E����=8a���W���N�P2Ip3�����"4��E=Zk,�@oTN���s����,`� 	f
 ��������y#�#��R�	X�|a2��X�6�A��3r��ct}<rC���dXK�d�u���6��0`���hn�Ю�\E��u!H��95�g���<�ʇ;z�H3ֽ݀��in�@���4A�ֱl� �l!P5M�r �ցa!¥]��	๋�
fk�)���d!f��C�!�0c7��b:�@��/Q���5��O"�4��FS��7A����Q�C��"�$/�z,e9�ۄ5�]���=3�n�q�8�<E�M���B;�*�*�Go%c5&��(�����!�E���]U9#��R��r>6�ht�!�9ee"y�I�����k5L�᭍	9��`Rz��ΐܡ�K[��`�$}�G�A��}_:~y�����|��g�9e�nH̷N	[�"�	����f��5�3y���Q�< �"��X��P�jи�L(��p{h�U:Ǧgk���#���/C����h���@��_7��ef� �o���p��kʉ�o,?Sq��X�m�L���F��yc�\�9�����/W'��R!��91���H}X۬�aU��NUu�ow�y�/�2��}bK�N�<DB���"���Mј�3�3�.v��(��d*��Ӊ�S_3ܷtG!ߐ�71�3�g����/���"}��D��Bi�
="�R�˸�a��E��E�e�X�ZF
�A�BA���4�	
��b��B*�=�lP���S��zⴾ�VLd�2L�Do*Z�`{_	��F<0�(�F�ýq�څX���У_;#8�J�n�z.��EL�X(�T��Q�r�0Lk�䈽�Q#Ǟ��d�J�V�#.*ȩ^#M8Sb�J��2�	r�F�A�MF���m�Ti�
0c�����q�HK��#���s��DuE���̔d��E�
��2(�$M�8B��A�!��G.1���U$A �Xa)��՝�ز��`B*�@�W����v�F`p�6�������?�"��[�4��P(75E�\���ǚW���PB�8>H;�X&!��E�/�4P�a���V1�(�щ�<������L�5��c]���Ё���2	�8�����<T3R�"�ǽ[�<0A�Y�e�@,�y{��qG
Z�"5�	1��Ү��PL$�KH-�Jb�S�%���IM�ZQa[��}�N��Y�=��8��x&����&�D̘t�K � �% R�L��X�@�!%�1#�M��-��q�n���D�m�o�&v�F���$�V3G!FK@"QMŰ��`#e��M��M4�F&�LJ��ێ���@��*��'�rr�6����R
I�CBw�������t�wsG��|I�MY���˞�7^`��Sf5/u
2��Ha�	7���2jnSBq�a`�(`a�
)�C[����PB�0�*-"�x���b�f}�Qൗ�f,����p���1F����B�zD�b���pH`�mD��E����A� �ڗ�->+���ɢ��$2ʽۃ��5Uӓ�P]R;�
s
�.���M����m��~�a����`T?(f&�;��	��K쁢�} �j9!@��	�T�Y����ʅ��hTB�ģ@⡊�xTǌnepuؘ�L���j�v[uė���	akBz���T����`=#ŐO��,=>eB��i
�ǁ[�0[�]���G<(dO�㧵Z����,z
���8������B��jѧ;a~<)_�i�h����9�Րt�$	09(����m<A��{s��� c9DLA��h����x�p���p3����W��,�#C���b���✼1�q����b����"ċ<c+M(��)z�DAhF!i����|�sǘ��Q�A��y�B��0Ljɑ�xƂ�0A����C���ET��Zĝ#��#CaQj"��+Sa\srP8�֦����,�2��^ȓ�#vv�c��Yl����k�(!Xℨ�ʂ99��n��#|�⻖�]+���dx4S��qk7SiB����ym�8�GQ���а�щ�ms�&)z��!Q�8D�A�:���O4�Da�<�キ�B;�Ĩ�S!d)P-�|��y�9����Vt��xb� �E#f��w�}с�qv��MbB���\��`��j�;'.0�m6I"� L᫂}c	"�hP�	�*L̲~Sg��fb�bC�U9_��n���!��g�PuKM!��&|�W�M
�C
ޫ��Ę��\�̳y�$�3�w�Y�Q�x�<$��ӡD�Ud� ��wTK���.g��j�3�	�
XC��"�[cp`F�p�Z4��"��Z�Gf�H���݇CYBMj�^�{a
:z�EM��;�hَ���ZV
"ۀ���x*W��w��l{	H=^�F�R�����҄]	��3�13-�=WTo�T��$!Bc�B����zp/!:)�b���i!��b]��h����"tk<�	�4֦c�"�!��r׆�]�^l���ŭ�s���*uZ�!�s��z�иiG��H!�,�PAdT�Qz���6��l#��/��F�It�Ã�EA��L\�f�!�-Yey�H��c���^�P����}=��C�=�"e�\1���"�ޯ]��0Ss}#Krf��k<f�5��T��wb7Ԟu7;�6\�
��u�>���ߚ��6���ƫ�BFU�Bꄊ9,� �����/���v�6���C*0�^y:f������!�;���[�ԕ=��+u��j�m�XQ���A���P�3��@�Ң�A	dO%%He!m$��i��"Fe�hΥ�܃n\,d�n�ǕGH�)���N� ��>F���&��؁P�k9r ���Yc�ÖU�s1gL5y�=�M��rEf&2U0$րSJ)�����z�1����(uW%��{�Ԗ����j�%��N0�D�:M�����t!Ǜ'c	�Ka�xJ\hYC�x�!�h!<V�X��}E�!#c�e&��0J�U�UR`��=�|Fp����B_�!N�(�mѰ��f�m��\x��q����u�UJ5�f�޽�ǵ����-A5��4_;'D��fh~g�{�G�n����@�b��I>���æ�8�Ep�r�n�����W	m��8
P�����7E� ������fi0���!�𲸁"�5�؜T�Z��vCi��
��ĬTbF���+rr�N ��l�������2��f�|��}��P�0�}u	PO�I��*(�کb�BB�ힿv<&�Ѯ��LX�|��K��wVw�?A�=�lAz4��
K���^*��G.U����S��'��Q}���ㅪŜm�]B�e.෫�K`/J��Z��/�A�}�ظ���5k*\A2�ܐ�#)d�29Y�3ض[�*L�@�#�C�D'�5�<J}	�W� �Vy@�Ta��C�9E�c(w������A�Pr�Ah�(E�NOv-0��B�H*�l�#6�d�m��ŘI����!$3<�F� ��
"���nO�:�<�{{jOT\�yn�+�|\�D��č-��htN���aDq��;��_ME0����8�@�ي�x.SF���B�SX���g�u�k����J!x�R�5s�x*Q�x�<+@S�a�kȱ�I#�������J���@�!���Y�]tri+��"���<��2��\���%Y�ѻ���0GΟX�C��<�_�7��O�A	�a��+n�Yy���}�q̾��D�a�h�;&V�8�a��o9TB����8���PB�4;U�\��)RJ���@� �K��4A�,>I�}<=9��<���{�<ˀ���h5b�o}�'p;/���U��^/l��-�n�'�uK�w�V+;����7q�.�p��S��1 p#b�(ȮtM�;5�/� �FW����׉��,��y��wd��{�$>�T�� `0�L0�M�8�����]4$�4GC+�An^<�q;&�&j:s9�4-�"LvmkZw�c��*,�+ �zL�K���y#1+�Ve)"K9���h�ѷ��h��B��Vq D�4Q��rG̊�.;�¡,	j�,�@V��ԁ���Qt�9P�f���&!b"ND�%��<BV���k�MA&2�W��U@��(i�A��ؔȇr�]�g*d̞gV܃$�[?>�ɏX��Z넉l��0[��d|`p�b����hz�O7��m�;w��s�	��n�츩7��aѻ�ı*E�vir��c�hJ��֎סb����^�:��f����3��d�C"���çu3�]0���3�9`��h�I$%e�X���*,�6CU!�]㙣�tPz�;'�Ie�Z�� ���1*ax��0Sh�����/)+RY��1�zsy�+4ڒz'��[tPBjC/E����	��" �	yUQ;�����s�,�GUKy�U֖M���&<�Z�\�0�� [�.�Hf�s����r�Wexכ���;~��&�詉��5M�����O!0w�Kw�n��x�4.x<@�4-���n�2��~Qƪ^�ۮ�Z��k*�M8��>�9�T���<��Wɮ�;��2)>d���$����r����@��3|�����[�
CG%���E�qN��h�uh�4���)GAC%�$"�"r6��͈IG��r��vws+�t���|;V��I2Q��̫�Z��[�k���$.��uǓf�������/�9�=*y�3��8���{�]�6�����8h2�eԺ�v���.�:x0�lU�j&��H�d$�_VB+����A��>����>�n��H a��.��;j�	�-\6�Na^�~3:g��
�AF���I-"���MC#68ni�(oq\�t�ϐ�cj?E�Q}��I�a��ة�y=~.���4�3�o�*���dbǃ
f�[_��y�Cy�<�(��i���		�zԁJ��,SA�x�TG�0J
���fX,j�X����0�.롾ř�zY���Dq�BZ�(�2�j �/Z@EAFDRAG���B�**�**%��"!x*!�*���0� ^]
�b�W�QdD�nUT�Z�Unܢ�uKՒ��������6piF�4�0�Ѕ��aY� �2"���+ ����5���Zm�Z��,7iߍ���x$�V�_�
P�=8����> ���E[ ���s�� L�c�鱤_��N)C5-&��=�ޯ�&Α��oqݓgA� wC����ݝg�$��>���|��Z�(�O�!�R�,�'n[������w���߈���Jn�����������C�Ï�~�=�N��@/5+�j$�GՇ#9�l;�#�/|��L� ��=:���dB�$F�@�l���F�}-���pn���Ö8�!3:^��8���l!s�`��z��a��3�B��٢��ټ 0���(�s`��)@�(B*�QHA�������V�@���d�)���N�����	��?��󊨎Х�]��M��uC� �W�)a���8����̄��t:pyr�߈	d�T7��׻h�?i���N��I	�����c�z�B�G�����M2�="�_V L!8�N.!�=�����5��X_8+��ߡ�Ѡ�o �H��0� Dc ��⇉�ڿ �˛���" ���6��be��<=/$6�Wxd�X��,��X���!�$LT���O9���@�]�)���$ r2��p8�bo�u��=�sV�%����)�m����aeƒ�N���`��X�-�}gVກ��%qK!�,X,Y�M$G��l�22L�l�+�cT$[7]k�;��o.-@f� !$Z >7�"�a�H=\�߫j�� Q�8��	��G��(u��&�����,{���v���)�����9�s��,�q�7Y��1�<����K��v)��7�=�!� �&j��s) of��6y��y �P%	;��>��@P������ۼ�?b��o��nD� M���1h� A����kp@���*��	u;Ó�z]�����ݞ��B�5ާ���ظ��(�A�d�tdp03�8$$��vV��I��S4 Q��}�'��p�H�"�%5Tǂ�v�q!{xS�/�R��k(a�Y_�����S�<z�G��m���K�1x�4�<`wxF�"��]�0�1Cf>��C�M����?X��_2`�f�M����~�f!��|"p8�˸=�y��$1I��6�CHq�*G�L��ǩ�h��7;�a&CiX;�C�2�q����ܑN$�T��