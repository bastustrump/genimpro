BZh91AY&SYZ��w�!_�rpg�����0����b8>                                       `  @  �   P ���@    
            �p � (      @    ' @    =�VR�� '�t�}�{����e&�t�	��C������zyx����=]�꙼�P����l��@���M�j��u�     ���s���\�<O{=.̜� NR�Gʞ�:ow���&��zhR�����詼j�-pGs���p�J/,�{0;)��t���@4@   �t      0 @K��ԥ�T�dG6Pxf�8�y�����=�٥^��)�U:s���:�a�i
^�5��s��]�S
�ޘ��]J�K��J�  U8ۛ(�;ro;�iI�Y.�����/!��u�Jޜ9N�y�^�E�{�U=�w�	.S���;"U'7;$^6�{<v�U�m���  Y     P  %�)^���u����W6���l�4�3/L���<O%�OVg6/{����=��н��8牔��=O d�W{�G���.�ZP   �  ��%c��jn< 9^��ҹg�^�R�4�6s����5��$���v#��Bx�OO*<�=���-y4�`�7e*�  
�9 �@ @ A�.�ȶnf^lPNlT绊/7�`����ʑ^^ ����oJ���{��6��͒U9�nwT�<� It(C6^=���媠    ��uR]s�r���< <�W�mnG�J���uDLL���^3*��� 9�+3^���ݛ�a�"��   �   = (  ` @h�rf����7w.��"���\��{��w���j�+CW���hr70g��Dzt��rw�i�d  {  N���6�G�����d�!�����T�c��{�y/!�p ���[����塹�,��@�                                 �  S�%)Q��d�=@ �d ��R�IT�@0�� d�@  	O(�LUU4�     &�I�@*�i�     L10�"��4�M�'���i��=454�A&�*R�&L�41 L�LMs�D���� �\zN�����w*"����UW���!@�@AS��(�b"G�����*܇�)���ţ���3�29��hhs��A9g���MXw�((��)���`AQx�pb�x���i �Q��3YC��"�
����y�������v��((��fCɇ�&��6l��s��Ϧ����m�������#�&Z��d��F�T���(����n�ᰄ&���f̓U��;K��1�-��q(�mXZ	eJU�U�`�̍�t*�w^I���j��5r���f�q9�U@� �ʌE�*쬫��vR�'��V�jM]�9��JBo���>á��縞lg��gJ�p���x��b��c�J����5Rn�����Q��}�Wc�.Օm�UU\����0R�D��[��z�+iMͳW)�R����I�FS��>S#,ڙx�Q�(�B�e�f�T�5�/-�J�EV�ꂼ�r^�X;7�b�I�u[�il�2�T��&���7�q
�R2�!;t��y3Q��a��Ŧ\n���nVܵ��伊̂��[��n�]�&}�C�a�x�y����7P@����%�;�xI#�*�s(f���꼏]CtsV�q�F$j��i�b+@�v�����8�kU̻p�@��$����)m���tjhf-&��A���I���W2���)���Ae���e^ڡ3�EkNV\����,�3�5U�l\5t�/L1^�����+��5�ꊖ�Q��]8e��r�;5�Ӥ�۬8��+�ec˸vf�F��!P��*&��m#vofL�͆�Vw&�z�'y$ګ�S.���a�2PXNÓ^����*�P��Vff\�W���V��M�,����إٺ�y{v���l�U����n�ӊ��S�ˬ��MP���a�&&�;������D]3W����˛��k6ì�.۪�n�n�յm�GZ��,5�]��_�9��-s=F�#Qv��h�z>��#wMԾq�5d܃+D���^�މY$b�m=�fb�Zv&�����-.�˩ �h�8�b�ʊ��uJfCaD��ʮ7nջ�☙��v�\�fu�6�\�To	�,�g�p��KR*B��y7uf_�*ݳw���Xyj,�2a������*SeM�f��d{�;x�e�;�EGr��ء�%h�0��˦s 4���՛�2syWgS5wz�Y���gȭD�;��
U5(.ÏT�,\8�+��x�u���̶�e�'i2��]u�n`x�hT�˗��[W,�S�)��J�O;�y��a�AX�p��2�1V�Q|��H̢��	b
QL%�VQ�PнJД�r��9VӔ(�t�QYF\9u���JʡzE�ݥ1��f��s	�Z��n��Z�ھ��W��e�4�Q�q3�On�+�n]������f���cZ�����S��)R☰^�)��P,�UElnxkeVɁ�nՌ�,H	Hw��(S�^�j+��Q��Fj�+Y�7��t5�U�5��,��J�2����yiT�;�T0v��ٴ\"���i�B$�ȡ�,�sl���X!�2�	SIĈc0�<�ެx,�oM3F���#���k�;�^"iD�c.��zd��te�l��*ͺ�j�-�F��a�&����cz�{	`d\ibB��[�Hb"�n���b�'J��K.3ux���cqV�R�ʶ텛�Ñ+��s44��MZ��7(��J�1Wj�V�M�m�p=/�Օ��=UWOn�
�kwwx�TӞ�o�U�SM�K2�QIb���V�.пM������l��b=;=A�9�V䳷A�7�8�F�V<69��	�/�V5ꏇC���V���s ��#Y~#/6��mZŊ�*�fma�DSVtQ �r,��J�K B-�{����vn]j��g[�ܽ\S0iU�Z�HS�ڬRU�!J1TFH���#KE��&R�\�!��б������;������V�Vm7��p���G�����$!{����$0S4�۪�,^�*����u,�ΰ�1vMf�6��t�'�YT������:HW�	�P�x�L��`y�����@a;.�L�.f�F�<�+^Ӽ�����x���e���6D��y�k)�v��a�E)u�Z���0v��V�R^�)̋�Lć���ecJ�&��֚�^�b�h<�	�v^7�C�%-��SU[D�wZQN��Qݢ��h��r��-��T�՗���yu^'7ۛ��{��J��T���&5yB�(EyL�dPWyWAǍX8m�uy(T��;4s�P<.no�uf��[t+3f�U1�6�d�U�6��2���~ת�ڤ�e���F�[n�z4Qĳ+r�jf*��J�i/�5�c.�խ�t�f�"�gu
��%���I��`�`���چ�[׀��zvB��M
�2T����b�"���g���*:1�jldqM��U8/[���3%ê=-t����[��6�ku��w��Z*,ViU+	e�B2�YV��s�F���q��l̠x���˺QV�I�Qħ���O_��6n����4�����R�"�Ἲ٭\�)��
���z���ձ�j�f�AӖ�M{�d[���w]�2վ�-A�"�hZ��̺O$P�vE&�
NRRnS��*!x���;j]Հ�w[��h��wK�8����X�K(g��X�	�v�]m��Z�*�Vy�h�ݚ�%�ÕG��ʫ�����;ahЫk`ҁ՘�PYw�Op���qnf5����l;j��
���o�uldV|Fj�`La�F�Jˇ�ֱ�B��n�˧�sv�`m�Vk��cA��[T��[b�'� ��{�e��:t�{�p���y�54^X���fNd�R��U��G{�MHڏf��WG(�WTEVV�2�������&L��Y���Q��Skk=�GpeYҦ0]���E)`�s�سbR���5���6�Ћ]����s^�Me�H{4&��Cn�f!��CkT����+Sm;Q%NdC�u�s3s2�v��©��!.[�r8��w����*i1T�٩�3��P��ں��lA!���V�Uv�F��6Q�wj�5�n׽Fݽ\p��)��X#F�"�:"6�0�*�$���\v.֭�Mf�/H����+t�dk����2㈼iDf��!ە�;	�.�u�Α��0�6E!"��N������qb�]��4)�6�@Ҧ��42\w�]3؃ᙗţ�(2�Xj���]I��[��T�*ޣ���mE.������3�ģ�EhH�7��(n���Y���	e�v6}�j����R�A����t	;[
�kNA;r�qڳmÔ�b��%���U�o���(
ݣ�������mb�۽ͣ~��v�i�<ݏ�K��;�5�d*��ƱS�y�B]��V͹L��ݲ��ih{�ϰ㣕CoNmS���ɹ�&I���Z7������!�w���]y�ti�R�:\U�pm��fl[�d*���Su����+XAU^�����0�̎a��;�zMU��g)׮M����;X�ڍ�R�L��ǚ�A�mT�m��Lm�k�ۦh�.���I]��c^�owcX����J����T���qT�Xu³U[��l=�՗/&�ދ��ޱ���Di�J+����+�(���?_[=yUQ��ͺ4�K2e2��[Ԏĕ�/H���;m��[*f���U�IU�׻�_�[6oe��HV�Z��N��չ4����R��36�kŐV�QXuX��+l���6"��lPt�Y�nf,����i���ױh��E�΅CQ��Y6�j�xV�#���/+�-4)=Q�:��r�v���ѯc��wIѬ�U����7yA!j�4Z��M���.�T�	��v��$��
�p^ځMgreԙ�)���c��\d��D}�R�Yb]ӳ���Wj��j�4�����ѱ1�F�0�A����˵t�
QK&RG*�d�m�#d�X��4n�ŅH��*��NfzE�nfK�6�:��וl�5jK�po�ݨ�]a�q�aǫ�v	G��늟�X��ȱ��,.���u�f��4`��Bc��̮��:��7k�fa��e�ԯ�ݭR��p.���n�N圪0C[�sf&��i�Ua;���P����:�,;qQ�ۚQķ�UGn�5Y0�*�d���)�5*�Kwlvn����a������M��Q ٳ��[6�o�K{k���Y�{0�1ǷR��7	9�=�*�7��qb� ��9�
!��y�v������[�U-���Υ��I�^4^�4��^�$��cn��p�b�6����+(�ŹV����g�3^�&a���6�����r�e��u��_�f۪U{Z�
!�t3) �e'�R��oY�8Bf����;��I��1�7�n�ņ��+��.ކ%U����q*�lw:��㧔'���+hԭ�/��<�U�b�1����c�v��髣YF�RۊX�J$�V�W4n�t��aO^-�ܒ��b�a��S������S�FΫW3"P����TZh[`��2m��(�S�6	���Z�IL�Z֐�ص�*�Cld9Mm����b�����.�t%�2�/j����4�wz.���n�KN�nG�:��"�Z��r���D�<��خ��U�������lFoqcb�af���I��wgwD�b�m��wM�nL�!�Ñ�n����j3(��of�ݛg�x�^����l�
(P�W�7e*M�X��e��BE����[n��
��e��L�P�jh�}�:����ֺ&��٪jU��uE(��5�ZTo.�,޹�iP����f�8,ɯmh;T2V^�zj�8YdRi��ī�*�(l�ʋ6��n^�۬�Ć�yC*b;]�	��5�x.U��OQ��i�T]�`/֝Q��#q�fbVV����K�+H�2�z�0�� �Ui��,�:×U)�R��P�����#�U)A����nj��e,��޺�7��Q��5�fa�0�<���m���7�-n��Vhn��WA뤠�5u�+m|���
{D`�9��
7�Uc���P�	U݋�*�Ʈ���v-�̗�[{{��u� �~��Dz �e�z�E�VZ�1���Zowõj-�.TUU�u����.�ܐ�#M]�n=�5kr���p�XHA���z���:����13��.�B=���$,J��a����AN�9�x�F���1�2�ɉ\a^�UWCe˚�tF,�ɉX&�f���ͳ	��2�jU��[�~�t��U#0�W��xꎻmۺ�l�f��Xl���R^e�.�˶o�]>��n���X�6c�̅[��/$�͟`���id"�̭�b�he��CHG9V������&�`l������-���y��Y���z^�ʡ�4#�
�,a��]ն0W�[��P|�1;nVU����;r�,onZ���fD��B���&e�z&cU��h����Ջ�C�qU��V(o�^ͷ��o.^��sow�����C��^����U׆x���6�a]�j�n'2:՛�u��mjV�rfeڒ��ϪVQ�4P�O2��#�5��n^�dnb����UY��ڸ�W��s�׋k2�~�}r�QͲm��t��ywB��۶�т�Ub�͗�Cy�2��b��F�e'�J�J��,T���������;���h*�T�P��޳��EF�%�����S���b�k��v��w�ufo]L�t�ە���.�OJ�fe�:w/V�-:f��ktE�d�H�q؛�h�����W&�{e�[�NB�V�K(�+�pố�KWk��Tm<�\猏�tշ���{�je�K�wQ8�0����3z9lnQ�t.��ZE,����)Խ�zX�FU�I��I�l���sDE!�Cyb�Gb�\�)W���4�2���WS��FWk	/Q��1he���U)���o�@�&�)Y�3��R�`�V�R&�n�U����1=�H^^k�03-�U��ve�n7v/tY;ǃT/������6�E�g��U�&�JE� Ͳ��:����b˾V7U[ۙ�w�����>ÎkK1yjf�2�.F�\��A:�f�c"7�7�C,6�d20Q�84f�e���̈D�a�K7+p�˸��QZ:mc͂T��I�#w�=V_��]ݡ��'�e�Yf��D9�㱵�ԬST���٧�b���G]F�]�t�´2\���i��UYz6��6K[�)m�*#
ӖNM��$u*۪�r��d�e3z^3E��[�{wu��ؔ�O6�_HY�!�,�����r��R~��Ua�/w�j��Ϥ�[j�st:�(])u����]]����6bfc՚����콬������[.� X[۩�\��F�C/hm)�zqG�!v;Q+{�Q�R�v�r�����/f�̎��"�bY�]���lVm���� �t��y�n�L�i��nM�ux2kp�\!a�b�%�n�\$T_akiu�,b�ٮ�T�U�,S��Y��<�b�$=���)���{5{6�I�3��oE���������^Д&⦆��t�q`\��sB#3los'��b��]	\��L�V���%�쭮��U��Rl�ڴ��F�i�0�^�%�U�S��^骣*��n�Jc�l��2M��+l6��J#3m�!`�b��ɢ��j��lb4feh:�Sx�]�F���lK�V����&R�k�oAV���錩�<�A��2ږ��������ffZ�&V�7N���Hf����Y�������3+%�(�Q˲�4^[Y�J\oI����0`Zz���f�3��jP+1��(,��I��wXYG���v��&���Ы�e�����i��wvu݋�}rK��X�����i�mǩT�����6m�˷�L3^l�����n��ٵZ��к���2�����DԗS�E@aZ��>�:G�0s�v��q�)�I�q�6�xЄ-�D�X/i�9�e��X�Ea�jȖ-άrd̵��47���7B�ӓ6���Qw�suɡT�^� Wv�(�v���E�p��h�K�
�ULƉ�oa[x���B�c�w��`�F�[,^�k/n�jR�n��dw����`�*M7�Z[EiF�]�f���i�FWm��6%��T���I����;�Й�k�c��J�<�Zn�[��C+s�F:,���gwLK���7֨��aJ�`����O
{rHʡoJUgF�¡U�NThLy���n�t��f��O�/sr����86ֹ��vJ�U4�X�:�UXU������9���L���ώ:���ώa���}���<����j��)��$��SN�^���]<�f��n��Q�mت��n�ޣc\�X�r�����ʜu1�6�W\i	1�瓊���/�ܡ�5y7Z\�簅v�ʹZ�rY��v�>9���^��[^	�s�<¾6��[st���d�tl��N:��� s�:N7=��G�Pu/�k<�M��B�����v�l�C�&)�m� ᇋ�*nO[q�ͺm7�3�����o�2sɬ�ݙ�:8�{k��D۞�i[�\f�Z&�9�d;X�g�]�'�LG��<�#���h^���l�L{�U/v�뗍ä����N�g���/%�U�I&���]W^yF��q�c˷c���4m$[.8S��h2u�����_9�Н�c\����d�z-!���b�y6����t��c�04�X����cB�I�Ξ��9�.���;�/c��r�۹fnݴ����s�N�6V�ƣ�7dԴn�5�#���A{A�l�N:z]q� �X�;<��;tmb��`By$��kp�)[�y���s�;;��N���g����躗�ݞD�3���xWt�����k��nڱ�'��y�^Ͷ��*ؗ�m�W:�L=:���{��[\��s�;�4uÆƶ�]�5�nh�ڞɗm���������֋b�z:�vy��+��Hs�{mS+2��L�l���9�cg�I��x�%�7��=�`�v޴G5v���Ƽ�U ;e0e8���V�Ef�Wd�Fy�zįV�m��4o;�5���Ff&'u����sOkd&]��9���=n��N:[ۖ���݊gg=d�wO\܋\�yokf\!ǫN�͝K���M�[������<��ʬ�W��R����K2�p�׳�x��i6��4�q��μ6v��K�=����5&��+t���q���p�:�4:�l�v�2���q��xr�_6�p��z�;T�݃n����glr�lY�6h���9�ggk�b�`k��i+=��8��F��6M�dn'6����jOi���k	�ﯠ��b�Ju���w��Ù��p�<��y�6�\:��bl�}N�{8�vɩ�ױ�k�J��<����G�4Cuswd�W�p"�X�n׳��!-=��\���g��y۳��]$s�;q������F1v���Eݻ{�{n#v��iM��q���[L������k������tiV�n'ہ9��W���<৶'��U��l�ps�u�t��&�n�Ƭf,8ݱh���.���9�q��k��Ѷ`�.5xv�ݳ�m�,�E�^rC�9\��z�t)ŷf5�3��"��7@�,������y6�mg�WkO	�,�n>3�go+��`ÇE���B&�"wr.���]ˈ�tY#�sV�/\����D�d�f8��[�s��|��������݆�[�<N[�8'��c�#���E���ޓ+j�Cs�ݎֲ�tR=_*'3�������^�d	=�bCmYZ�n� mu�mϮ��-�:gn+I�T�m�A�n1�,ݍl�Nљ��������i��z�pvSe,gk�gc�ۤ������Z�ꛅ��qy͋��'�~x��V�<뎲��qm��<�Z�����RV&�Ѷ,2���6;+�9��i;��\�Kۗ�ɕ�"����fwrDۆ�aF^�r�˩ۈ4��m��&�R�&�9��+�����ְ��'/sr��h;�;lukЪ���7g�ݼ��OHM�8Pu�2C`�N�ܬ�^�� ���nӷ)��������e��2�d㘺���n7Q�v�ⳤ�Ͷ���݈uʪ�m��\un�cߥ�|��պ͸�^{W�8��cx�x�l]���x٢��Z�laܧS��v���y$�ֆ7�����Yח�hR�P�]7/k�oM���GX�����z紷.���=�Oj�hs�vX�sGk�
.�n�1����ll+���yy{y�g����<kk.v��qz��+{[׫��X���rwq'����.���9�p薺q�ׯd�m�W,�A��d�Ɨ�t�ؘ�[)�1����n��l���P[��o�����髫fWp��v��:��w����v�|��<��ն�I��]�s����@�fY�[q���v{uѻ+�Ƕވ�=���ZӶ*:���A�c�u��;�;fu��C����)*��&om<� �%�ՔW�$��@�i�]�5!�B;�n�6��r�l���������lv����R���:��#ۙ�><7�sv�!=3�lT��j�;�Kzq�.yݼ�s��녖����k�#q+ύ�f��N�n�4�[�Ѱ��4���7T{�j���x��IF;��[6� �lq���mțG.
w�qJ���6kc,D^;l�y����Ҟ!���ʶ9�'v�í��w݌�9��m�wi�&����E9�ƺ�2���'dv��v�uZG����zU9Y�=Cme�*Vd��q��˜��-v�C5U�W)�s���s픴<�K�Z��{��pp�c����:T�(�n��E�c�ӗc]v��GOquY,���V�o�7��α��i8����$��e�}�?|w��v���n<�f��8N�u۬g��6c���݇��@�Gc��>����<�i�'���8�i��`�ق�X:C�F��9�Q2�m�l<��m�sǳ���ǧ4�����0������n���1�g���W��ܜ��Ks�����g�s�^7<;�n�1��ۛq����nM[nn��|ҝ���zX�uΘ��s�7���jw��97$	��vtn	���j|���l�X�����O>��q�����+�e���o7n[�{w;πv;7���)����v�q�h�c�۲ؑ�ܖ1t<q��EG��jZ;�w8�%�n�'n��`1��&Getb���c���GC$oP����Ǵ[��g�Lyy�C���&7�&nt<]:8� ��鮍���M��`-�I7�:f,�:�t�]���I�ۏbB�N�]7�wq���6���.�d���{Yݘ�ͤ�E�ᱮ^Cgq��M��n��oS�}�*�96n�V�Ս�d6��6�v����|��Fv坻��z�G%���]��D�:��ȋ�s[zC��L#��9�a�Ǘ������L'r#6�\t.ɹY�m�7��-�)s�=��y\�������mRv���w��ۯ�y�G���P8��݉1�1c��dP^�FM�1�qۭ�\��v�=Z{,n��gvt�۶��]OF�<�O[�7Z(�T���������\��ͨ�7S�����G-��J����v�^������'V����|���������g<5[B�j��(飃��Ɍ�n�e�Qw��.��f3GlCFv{mc>��F�wBݧ㇍�=�Mq���!���և���1�]SNyCӻ�\vG;���g���ֵv���Թwk�;[&��N����;9��;�]r��ņ��v�L�27lh�O�I���Ov�<�z�\�����z�R�ٚ{a�˰
���y�o8\�	٬�������7��&�9]�p�u��qk�#��p�)v�aƚ�G��wWA����q��Ғ�١��ۨ�%ٻg���7k�
�󜌺]�4&�W.��[��uZg/1�J8y��q4<-�H��͎qź�m�3��bN���ڭ؝vL�\v+y���.Wpu�񇎮�<�q�C���s��h�v��;�dleL��اs���n@�7����cc�ls����͎�����y��\Mgs��mi�ƪ�v��w�3��)�s�;iz�9-{lJ��l�\��ћg�Q���Oc�g<���Uڧl�p.�s�-�Ȼ�3��v����
tfns�� /cT���=�� ��4"��G�P�x���!�sی�F���������i;g6)X�p*��d}��'�k����um�6�ukYkx�n8�=Q�Xヷ1g=���n����N�8�n�c�0V"�9��P�c�OK��K�:Ǔ�n����Xm�ȃ���v�}����V9���&�Ԋ:i&�)k�t��z����;[ۭ��z;V,v�+�$8O��5v7�iwUa�\q���Inz���FW�������{w�ιlu�0Hc�|Џ���s�G����'2�#�k��;��:ܽq��OZ7~���]mq���H�c(%����B!q�A���ɠƍ�b������k�Lm�v��qո��[�&�N(4۶�W]�/�C�'&���.�vnqI[l�4\��vi������s�v�sv�ܘ���m,:#6��c�u�q\sK�np��m-�s�]��	�����c��W�璺�f�0�u�HM�mt����6�7bq�u=��Je6m���!���u��rsƶ��y����#ں�)��<�ώ<=Gv�c5k��a�qN�n��[;�d�І��Lܞ�rZ�뢼(j������n:3n=�ݹ�t�_I���{���iܷF8���η]�-@a{(��3����5O�d��XK�Gm�Ã��n�Y6�3��ucE��u9{B<.+u��i�r�j�qχ�/����3Ή��q�Y�-��F�˫��.�.� ��'�ن�k&����]�{Z�utO9�[��[���rxkk]��=�n���F���zM�R6۴�;8����@דj�g.r�7���ڗ�y�T3/m�t���.ڹ�s=c�G=�{]����T��.�v�l�
��r#�xe�z�,��Vy�p��2}�~��m�p>�[+�:x�<m�ݑ����*���1�uxXKy�F�:w��!{:�y��Q�u�v�l�m�+�7Y�-�/���vm�t�F(nl�6���g�,tskO.�Lg��cN�m9{	�W�Kse��:�Jm���9��Cö��y�7��e��9�&�ƈ�x+�۴w8�N�.3�C�n{uw�{{n�����a��$���-s�p}��"�-l9}������:��6d�<��i�?�z|�̓�������*_��['�<��s��M̺�,�f]�_/dΥ��7���C*vY��R3�^&�����Z.�L5a[^M�!��� ���r4�uv���{�:#��xۭ�wGr$�F�Ń=�<�����b|b-c!Xڱ�����gڢ]�o �:f[yW�ḁʫ'=�ڡ������ܭ�VB��4����Ӄ���Z�va�`yId܅E����d�ͥ@��S�k�:�8KFWWQޮÛ�G�av$Q6w}��4л2�VdW��J��}ø�mN��1�J��2�5���%:��ڵ�u�C�+W�mS���C�*jĢOe��GV�L��}y؞8;,87�f�k�>������ ��3��%��࠴{�x
���������Ѡ�E���ui�3n͇����x�S�$��xv����]�r��7.m��K�o�]{:�{v��u�i��Mq�Z2C�i���
 xz�o�����e�e<��{����3*�����Q��xxϹ�Z����ʩy-踰(#YY��*])��C �fb��؆NB�1v�j]Ҽ�v�[5N8�U�/�屷���Ӏ��-�y����r�Ѥ�%����"j��2�l�;E����$��W#��n�����64�]vVN	Z�[B6�^C��xRJ5�2���̍k�q��&�Gq�hL��9:�������\{��S3-�D�����3����+�e��xx�Q�h��N0��:����h�w�X�B�u[[��ްэ�`ێ�n�K$��kYR�T���� {�Y�����ֳ�f��J�` r����s��u�n�����ک���Vsd��� ��R�5��!5kxS5��^k�Zl�P"�^8��w�����ۡ��n�h�����9�u�7��Ԋ����V+4ZU[���j��i�xen�}.�5�gU���ٺX���m�hfɪڹt��U���z$=�o:�Ś7n*'cA�ٌb�q�]�����d8��sKX^����P�k*\�v�����BeVM�e����ʸ�ށ9`x{�;{�����V`�G��<vo��w�7(U5����)� �0K�n�
^�
��M�� ��w8��]�-hJ#F�ˏ�q��2������"\�[[n�����;���2MRλ�Y��ӗC�)�i��h;S8f+&r�=�up[��Mpέ3�S��z��/n�έ\��j��I-+��c�!��-H`�B��pw{7P��"ε�A))����Vи&;�Y�b�ӷ*��1m�{O)�H���%u�fJw+!Ow���u${ye���Q�T�f��1ٖ	�aV���_u�ս룩)�e-s�����i����uh���:�A�v���P\Iu���U��?EYW�t'��{��<3�ᚯ��Q�< UJV��v2�pP�����s{dֲ�kx �ԕ_-5�b8.�\��Z^Adɱ���i��� �B��gpoP�J�V����C�m�XN���w���B˼7�	3�R�zb��}Z7�19�P9��Ub��/�6�:���e7u}�1���b�Mu�ճa�w/T�wKZG77c�W^�8f���r�.��[��vfmRʬ����G-q{��ʝ6��#���z�d��ֶN�T��m9���mm���73Lk��7�-��sǝ�nˮ}����tXi��%�uU���/d�D���vMχ���u���1�L�SmH��^ ,@��-�of�&U��{�m)Y�vy��n���,�(i��X.�4ý�<�uc��[�h�N�OU����c�CU^�a�������o3r�P�T��\���yR�:ЗT�fS��C���kz([WH�I��s�9}���o��l�}E�R���[������C*�����R�O���U�Zט�s"�CQ��_UN�u������ȴ����e��专ٸ�����o#�O;�[��~��*�Bu1��u�b�v��&^�Xv5XP�8�V�.�9ZY�1�7)�ޤ)�9�[��nև�Elb�(�[���k�Y��x�m���
��T:]^����`�N��Ye�d%��@xb�m�d� �'' ������hv+F�ʱ��LK(~4�qBpɻ��5�[��x�Lk�}d�	ى^��"`�V��>�M����FY9]�������v;�x�w0�L������������c0j�:��{�0�oo��=��/f��BA��[�v1z�p��ʕ�ۅ���X�ᇷ&�wy�Dn;�ӭ��v�T�������֬t\�Uա�b��3�M�W����T�V�j��s2Cn��9Ԃ�ޠ�.����JX'��z5�}�-���n���Ԋ�����|zo%����ƗWi��ܪ���u���U��&��%Ӭ�׶�R�<�X���[t+)>��x��Ō��dK;3���{ޫ�pG�Y�W���Oq]��� 5�f�eh<��gH..�,���x
��ڹ��5�p�Y�>��)����U����|:��eJ"^��z�kd�:c����[�s*��P�W[	���Y��_7h�t�ݱ7R%�Ԋ�Z�'�;�`�k���0��|�IjUY�����uLO6��ee������X���z���<qYëX�lcZȆ�q{1�ٜ�n�L��W�G]�Jf�
���$t���[��lTѵP��nZ&M]�S��U�wZ�jN^����{X���;�bL��]zv���O��5n���t����/P�����͵
:{i���wuw#�ړi�eש��,���a�v�^��aLV[�T��8%�3��7�q"����h����koh�/mX�u�Gk+��;�)L ���X$����{g^�!p��ڦv���n����c껝6�&�}K6�oѽp�:ѕ�`��On�C�˲�&>�eާc����i+6�kevڭ�T�M���g��쇤��Yy��J�������<3Q�fːƍ,)��1�W��z�m�����
R�"��#,�n�*v������@�ڗ2dF·�je�쀭uFCg��n�p�wB�wN��n�c:��k�n���+v���2l}S�������ݴ�Îz�r���v�K�6�*]�u'��a�m�7{j�ù�OZו\�u���.�2�*�Yܪ�E֥�kx
�)��:gZg�������DU�I#����x!���^��p����d�7H��/qJ�$Td��K�r�_ڏk���SEV��^�ۯ6��L7��W ���~�����������/K�ֹ�5�Fw�F�dA� �0]\��+��N�;�M�˳�ۧ��їm��;����u�W=����c]X[�w
є�n��8�:�'�y;�����[�]�7h8���o[�܊�Sq�խ�:M���lkcl���+v��A�BN�!��&�ֶ烠=�&�^�Y����g�q���r�{��2���ؼ$�S;��N���[��溇�)��NK�/�n�'E(�jE\���vu״������e� T����dэ�;[۶�׎�=s�=�i���]�cj��.��������qϥ�h`ݻ>#�ڝ�����{'F���9��9��Wc�KZ�w�b��qdU�rn9^�v�G����[)�oh��n}�5{X�9ԥ���u��<�$��x.�����Z]ӃG	������c�����=z��V8�y���y^we��=��m�g=h��q�b<�;Kv{�ny��g9����v�/#�޶�̇j;s��b��.{[B��s�z��ٕ��:��ENyr;Q:6�[k�o6ݸ�6���j�웷U�r�;�3]b/8|ɽm�Ӎ�<k������8�q�e�ݰ��.n����.Ǎ��l��GP�3�g2nɓ��n��v����m�^�@\'süF�n�k�.��G�{^�%��.�v^ۢ̔�c��u����{#��t��p�5;�oغ�P��6{#��N�e5k=�v۴W昂���7=?m����y���	����x�(���t���=��a熳�뒆����(c���h	����Η��g���b�i��t�d���٭���07mR'v�[�u�Rs=�y� q�hg��%�N�ݫ�x!�u�uY�������^:G�sMF��y�v�q�p�fDGJ�{gu�)����8;g�>�5��Ě��]0Q��2�.N{A/�sv���ݽ�M����I�H��-�C�C�Z��Ec3)3���D�����	��XSM1�����"z�B(9[�cs�n���V�J��w��{�xx$P  L�
��e��WJ�e��y��{����C��|��{p^���{�Y��x���{�ti��;Ā�H@�v� ��� e3U 7�fHN[��<=�u�� >Lk�,���i��	3K�s������ϵ��@��0�&n����ƪ�=�Y 滌HI�g�t�W|�sW��)�}���c��=���I�@�P g۰	0n��`$����[�]�L��޸�%�{����!}�@7��I<��h\�0�D���U�=,*�4&WG� ���wƠ��B�����n����e��HI$#�  z�܀B��.�l�bB_;��k��n&3~ᖻ� �k�Ԓ�I�s�� d�� xa�� �l#6�'f��ٍ/���Z�V߱���M�]�[��NvާNJ����HnA��:���E�ۢ;���G�::2),`T���ӵ��(��㊱���d3];��]��oa`S<1n]�A�]S�T�;#�Xۥ۶��cO\�79�p�r���N�jƶ�OY�5&ö�l�l�Q%K[<k������=x�� �`�K���8�n�O!�d��<��7vyp�m��7Vrywn�6�8ڜV�>�uɱ�߂'������u�}��M���y���z���Q�����|�؎�$����ƛ����Z�3�Nv�.\=���>����L��H�o����#(�Q�P���!��z#^bm��5��Ư+_6dy�UE ���C���A�5�����o_:�Wt�H�PD�8�=֚kه�ASI!Ӻ;���k����ޫ�z���YF6�PIgA�}��Z�������n��7��X�PD�g�s����v��ē��2$��� ax�=�J��.��䮅���R>6���rQT]͹bF��{��~�����U�1�;����;�un��z�%t��4q���a�#
(�m�-�lApU�$��̂ʄ�f��b���0nb^x �y���y:!�h!�To� �b���x?�����%"O}������<�wä㉱>F«��!4�(���YD�kI=�bh�e	dw������f�{����h�f

J�"1`��h�`56�r�b��,�ňT=�(�$deU:5
�77�z�b�����Cr*�u��Cq�	!D�F0]���p���+��8�v�UQ�X*�$�#Bo.3!��L޻ݱ�<A(�QqA��APL�\QK��(��ED�?��~P�H�j2n��V8=tku�O]�vlfH�3���M�&R���_�?���_��T�WH4E1�xrr���K�Yttk�taw�W�Nf�"�	l��8Y�c�#��Ac��"��B�X�x5W�9	��	H�F�n�Hv�g�I����c�ŦGvs������j� F������k�!JR��E�=�K(���߯8��I��M��ea�(R�c���������4����)	�³k�M8b�i5��×E�X9���"1�/�	Sr�8lCzne�-Y�y�,:&�.0�!Ȑ��N�B�c��I(
((��j�8vm�;�8��r�*,�G,��o���&�Z�eoigN�*�t�T�VU����C׊@^(1c�P�ߝ��}gr��0�-��psB����{+��~;{^Nh�A��=��:h_4�4̊$�6v�n�3�&�w��k�1�_oz��a����Dd���b��<�EHx�k�i�����t0�Y�{��t+���I�mH$e���4x�������b���z=x���|��Vq��,Z����\G	��ƈ���D�(�T�UfW����e�=w*���7=�����K���Oٞ�++N���7���V�Ky����v�}/��z}�k��I��^/��U�����IE�H/qU����5u��|
�,k
�$�IW�� ���G8m�(��-��6�R78�\�`-n�Ƹ\��\�t�7X��u�݂x�ѷ&��Rx�舜)���#$pZ>�k��w�3V-���b�qӠ�����XN@�*�M���/7i�,g�\�����,��k~'=�u�x>��p0q�W����7v��]�l�A�����U�4�w�߼ _o$>~պ���δ�Gm��3CF�D�]���]�pK�΃7tYɅ�C��p�|MA�!F$r'#
ŝ��6Qݪ�
EP�.�{�{�֯��wP,������Ә��+��:CE �'Ȅn�|J);.
>i��	LU�s�as��7\{q�\��:q=s��W�78*1�M��:r�z�E��vNݴ#՗��o<*����v޲ݽ���x���z�����lܷ��d�����.��<���q��:5{q�&�����5,�r��9�i#���99۵���M�\���z|G���Nt�i:P��ں��]�:�v�$	&�p���BQ{���Gm]e�m��g�4�N^Vh���Y�gi\ݻ�����J��욷<ޖpֻ��P�����sͱ�S��_[�)#
yOl;��"��&ӂ ���V��|��#֖BR�O���}bmT�i���gӞ�a�XR(T��)H�uC��> �I\k:/J�d��cU���>!2Xm) )�ݒ�/1��MQE���y���|=�V����W%Dh�5e��=�Gu]�x�����3���}�\���/~$�V� >fn�O+_�ρ@�Y.F��"�CX:��/�ך�E�\�Ie&�LH����0����Ch,�7��Q;kD�Y}� ��.P/�K��U��!�=��kfێ@��a��Nk6�'�q.�߭||'�lC�U�Ŷ�7����J��rh�׫;��'ڬ_ޘb���ai�C>����c��}S�Y%�)@�:ó�S�'�j�%�B4`�մ���":���䉾/������0����jVc��=�����崸b�8J�������/<H ���xx/+�è��p뽏ZM��)FFp#�ő]���|��X�I�����m�Ԏ�NB"s�n.g�+�X�O}��2��"7>�c��5b
�FN�&�nB�q�\�_j�^R�RL$������3.��˻D�{j�52=���*'���%������o�u���Ϛ�ή��K<��y�U>�e����ێxY5�l&�tB�wٽN:�&�G���`X�Wb��"m�<��u.�Ssэ�h����i�Tm|<<>����j��[�e��ۿ6���!3��>	#�$��|3�D�#8�h'J{�>��wõ7�-�� �s�n9"㌓1���-��L���b�]��%eEUQ�qq�F���U���U**7aoz�7�.��zWYx��_<ť�Y��n��t(\��Z�ƚ���;F�]��`��X"����3�i��S�(�/�3�J�R�Hr�[�I��EAH��2� �!�g�p��tc9ޘ�]ً��w�d��PuPE�b��!r�aJl�!)��:I�(:��*BU7��7����-b�����	���{�y��zls�5:�O���j�k�����^���E�ȠA9�M�uxl7�`�ŷ���S;�.�`ЬP
@A{��9¾xU���Z����ZCh}�<>|�?�&Ir�e2���r�o]��J�"�b�@S�����O3VF�<�E����$��PnF�Q���`���m���Pʘ	�}�� *��ƅo��
�q��nnP��@p]��=�>�$hS1|l^� 4��M
�&*9Ya�D���ɒAE�Yo��{��f>:���.���5�h�wR�z�q��²l�ơ�5��Y0��*��U|��d��)!.x�F�1K{��:d�j���;b�`6��|'��8�1�,��ʒj*ϛ�m����%�]�[����)//&�f��t.̅4�b)I$�"�h@ܝ�Jlβv��U�T'J��ä�<2�L�b�1m�[�&b3
۪�6g��=�T�Y��Q!�W����k��W��� ���%8 ��qH[^�}�}_��'�\~T2������L�B�e���h��%��H��jcc�$>�����jQ��'��*�*))3#�$Q`��檫	I#R���z5�k���M8��F}��Em�8�8�S�xx�|Gӂ�A�	=�|����K���XT����������xw�˻-j�0��s^�AMYބ{w&=']��]Ge�����p�'6+s4����}[�l\uog������y��ۘ:�q�'9u�qTOn�E��v�]%跢�Wz�	�v�y��;�t��N��W8ݵdu5m��W�x�۞{&t�Ob��ki�{M���<�n�	�5ֻ.��=����>+�Q�j��:D�^�⳱s`�#�SMqb'�B ���&�I��~m�����us��;�:���ܡm�����K����_s��N���:���dP��E�rW5b��]�ӻ�iD����v�7z\)�
@�r#�����I�>�p\���vbC�g9��Ag���_=��ӏ�djP7�鮗�ݦ2*.j�T{ޖaB�zI=m����NW�xg5�����! +~���J(�h�`I0������i��Q�h`��$W�!{�U���K�=�C�!�ޯ�r$� �2I�>�����=_:�hh����]�$d�M^~mk�:�2
,R*�#:o�g%_vd߹�-'!���(�&���_� xb�&���筡�b�I
��{=�[����xu���r��_k3���9�M�vK�=�bK�v�YnZYhQ�ϒ�,/��2����n�nb%4m�RPt!&.)$j#4
I"�xh�pL��4��)6YCQ-�"�I0���8�SM4D �(�T��L���
��{��|����"h M�٣N�䲁�g��u��/.KÇf�\9S~�A�Q�z�Bo��$�⌘$1ȍ�����n�/x=���mߚ�sm��ttl��M�B�g�G��?B��ߛ�w/���0$�	$Bs!�q
=�,;1G��$S"ab����EQF*���=�U�kGD��܌�#)5�\N����2Uǹ/���w����&ӛ���H{����3�=Ϸ��M���U�kO8��.䧋.Ź��1�Гس'[����-�@M�$Q�#(o�B��<I�xp�z_'�ȇ�@8-ݡ��ФP6PJ@dq!��{�D��E��|�m#��1`_���}�x
�}�^֞�#D��O��e��7�}� ~��8:�G�<��?����A9�ک�e�)���ڬI:O����M�o��λ�/�"��RwwF�`�<ҥ���M�wDݲ�5D��3+7V� b��a(zL���ש
-�|�u}�:nr�Vo�?')�s����SN�}��sM��2�;�i�_�YYד�S�q��Q^>믜��g���D{rB��]Ѳ�uҢ��ɸ�d��J�hLb�g,P-���7C�\��4Ea7�z��^�
ʖK"�L���Su��d?U�9����[D�[��`XԊDJL��$K5B�aҩ�;��Ifф}z�.�=�4f��Tc7D�`p Zr	B�䌡N@	��Xi?��<1Z�~�^d(l���5��R�tTpZM��es^hÂ��3	X0,J�f+�p����.��3��ly�Vl�]�J}!�R���b�"�О9*�d�Ob8�k_��~;{�Q!�34�sc���j�!���lJ�e����7{j����LH�&S��],��l1Q"�@i-P$�W�P�Y�����0M�`B4HD�Ԇ��R����0�Y��8�mN+6�t�ek�ί��nY�^+�픒[�PuXR
f��نO!�C±�c���x6b�ʹV�mξ��ZW}�A"�M���m ȣ� ��Yp���*������F:�uT�G�
4|����.6�����uE��UV��������0�]�_+�-����7�.����w?X��A��!\�Zr�^NR�<���Ԅ��p<�0mvL�P62��ݨ^�q\b%��>�u���7����콂�OF�������Ėw[�؁����Kc�(�"���8^�]�é�ˎ42(Z
V��!}�͵�e�y;T��k���#M����{+EWIQ���,���Y����x�� X4s҈ְ��wguf�v���4��7/���[]�����R&(e�2��������Ơ���ݜ�I]�pXzu�������-�K�VPv7:��)/��6�׎=OiJ��O���
��_D�E��>��?!b�ȜO��\��&��a�P�����H@8���p!zB]�0�@�*7]���)9�ł�EF�>��Zë2!N؅�5�e��O������o�����0����6�&���'�%�X�M�Fm2&����x$+���)*6jk�)�>���MO�#}�W��ww�ۍ�b��9磬]�������W�ulBH]�����6"��CqFș�#�Y�������}!�z�U�[:������v��u1�e�����eY�x�H�1�Q{s<����]����*\T�߈����~�l��R���V��6�M��'���'ڣ�Н�������3�$a�|,�э�c�����
gD�>�
��>�M!�W{�ı���*�.�\�šc4����w����G�|~�F�,8 r5^������c if�H�A�!��26��0؇ē#l5I"�J�wx���L&�}��!�����F#~���@��*S�2b�J$Q���"�B�� �ׇ��w����F���ݻ��b�P�n�.���3 e���}� J�f?������+��۫1uM&g�2��}���[��No��q��!�� M¾���`8ˌ�wǸ�B�o�?�� m�k�\wE�mXgm�%:h�2@s��n�]�Xd���Ͽ�=���"�ưc	mV.�| [�	�9���6!�n��T0��a�o6��s[��J�����E%׎��Y�k/}9�N?�/�c�t����3-o��8f�k4���^ 0y�z!ƻߪ�M!N��X8�hᜳ'�0���q��X�3fTw���{���i�_UXz&Y�sT2����a\�W�H�Bm
�z�& �~�@�t�&����5�W�"��� ��*��.���X�^R�����SH-�{�l�OFu���Pai=/��$&����=����M��M�"QD��~^h:�����Κ��}u�d�hQ ��&,O�]Y�82�]w���Lp�0{T"".NX��?�ݖh�YEffC����&F���vp��1��ϒ@"A$}*<�2�<w;�N��d�dɪ\-�\kx��9�2@H�'{Mq���Wn-�����(��ݎy�U�箶u�hmY����=�O`���۝J�u�B�sٵ�nv�8/]�7���=�<�I�Woir���+v�p9�k�S�ί@�s&K�')�;%�����
����&5���;��eݧ&��v��z8�Q�;=���F�⇪�m��W��.G�	����'ju���ͭY�"�L�(ӹŎM�Im�]�U�x���׺v-�H2�=�"��Ӊ�-2�L�j���n�}��ѫ����0H�QO�))IR0.<)��[���*�n4?�Ͽ�����h?�����03�ڷ��Xr����P���"ّ:��Lр�g�����$m�$FE�8�}��=<A��{�2�5A���ܺ���Z}�á�utf�M�5�V)@b_�i�^���%�A��)�Y>"�@�қ���|�,��溩��A5��攰�ٚ��N����˚�`��A�GT��#�=ĕ�⪎Sd�eR"���f5RYHNNR^�]d�E\K�����������!��"�ׂ��w��e�B��G��|u�"X6h� ��q���m�!ԝ���(CO����0��>�z>�J�i�en��9�����I��9p����>P�9��V˻��+�U�n�ZqX�M@V�y���-�Wl�� �P�`��>T����T$�������vD�_�b���``r��
�DJ��T�"� �#a��-c��OՈe4�w:���C,��g/��q��YUx�j�30��߈D�<i!=�����i�o�U���P���ArX)�t�!�3�{�����4~���F,:!��\��D�ϠT�{�I/�@ݿJ��_�b9*B��/G���x���Q�q'�����u0'�֯���}������=�y]75�2,V�"����>o��9�����qT�EY�&��=54��E����ڪ��Lw�5TC,�J�z�`�)��M��0<:Ci�y���ϯuE�-1�n뭓�I�H�"��3�Aߋ�&�;rpB����M]�Ջe�:�.�q�dNsU��= !l݌�~���O6��n�gf�����Ð�ޱyx�vN����k7m ~�|1m�icRAb&�m���H}�U�a�hL�kn��\�)
�I(�g�f�}Tb�b�ԳtE��o	<é42s�ϕ�b��.�x�\
fpO�������NW.`L�w^��	��Q�f��q�BSHzCS�ϽU�/}Ż�$��+~��V�
6r̆��;7�S�����ܢ{x�~k��� G�TE���%
G!eD��ݴ4QH+KT�{��g��Mkyn�ɸ��e�][׼x�����@��@�Į����6Ƞ>�j�Lj��E�C���45��]?Z]����ﾮx��y_<��0X6,Q��cB����{J��e�w\o̶|A���t���2��c�ڣ��de�s��%��p�e7^D�� �xȊ*�X�ﮰlI-�x{�gE��sc0������`[ψT��u����������f܉E
�D�L7�=���9��a�*�z�mdBF�f	)(1�R��l���m�\��be�{A����A�L�DTXRO�i���7��b����E�8Ѯ}Tbu	�8^�}��W;�]��uט}L���da�k��``I�g�x(�O �Ϻ��0��2�on���)�=�����"A��j���~�la��~����8�"w�)s�%QQ�2
" �i�c�jG{��hd�:!F(��wg�1(���ۯ]H,�:Ç�WJ�V$�n�B����+�� <�� Xɤ���	���H,���߮�O2͌�� a9�Ìv����W�N�_[�P���n���N�D��{������`pd�T�'h���貱�a�+M����VI����2}����Y=��rCi24�ݵ~	����?T^��0�=�|p��S���[!؉DzM��\�Ӊ�m���-@GK�qӬ���:^v�i���G�3�8��߿y˾�DJH6P�4@"�,:�Ĕ��w׀�u%�����X+X�&�
D��n���ɗ���
ݸ2���Z��d��Ii+��������`��} �ld�Ї�֛ ���Ըl@�?�~;�����A<�.��?��&�W����b�)��W1l8���� )4�++'�kܺ����wW��34Ȓ�����L$�;��w��fY~�_���q8Q���{}��mz����nn� �%3l��x����Ͱ�c�O��h�þ��=-EDA��b�=��_��=�It��Y���te�r���m&�`�0g�w��Y�
H�{U�&Xm�d�r�� �{�"U+kE(*��	Tsj�杞W�E��'4��Yh)�.�#ww��R�Q��=W�7|E*b��u�r�UQs&Ų��.=1#׮�W�Y�n����V���1����ǖ0Wf��M�K��%�\�������[]l��lu�c�v��s��m�3ն�8Hw��!-�9�{��$����ͳ�p�vA��:v�u��6�OU!�	r�1֓���筩��s��{O@m�ut&2gk�6Pvd�#gn�E����nsb2N3gp���W�|=n��|)%�m�����l�m;d�q����L4RDA*M9�"����L�͹'��볖�`��֜ӳ}�s���x��vA&v����E���8��|���w�{_<�y��1�g������F�z�˼]~�g�	G�C��DE�����#$���Q�i�@��fu��I���:a�?pl0��!��>~>�l���U�0�v�g�-$;öK�ְRĚ1 ��#u*�����}�	@�#�yX��ĘhHo�bB�?9̜~�$�>��/�i�I���H�xp>�� ~�*�pm40-�Z�7A0$��X�"�PGTV+��ʭ��f���@��H%I����C����`��BM	+8\{/��i�t�ik�w��"q'��.����`��ru�lHm%s�U���v��ڟ1
g-��'P� y�W���u�G�)!�ImP�� �N�]��3DRC�%��_V�T��dHa�"L$��&
O <��ࡓhta���/щ�+.U0E��₊�z�f�[���������B�{M�֎�Y�m��3ǳ����v���xݻE��G���xQ���@�,�}�I��C��X-��lB���S�C��8s�P-�^����Q����~�wpm�۵�y��������w�K�$��A���\Jrh��,�\\���],M���s�N���g�}���9�O�K�9����ϞW=L ��h:���k����3�����J�x-bR;q`q$��[!F���Q�&�7�����>���1k��X��jʺI�a�C'�X��=+�B`L��-_��� �FQT��m�Q@�un2��$��ɒ���)YG�}�_8b�S�L2Fg]��!Ć���"jIA�����0G�{� ({k�7�V_�'���!�}�^-�c �-����r?f�������-׀�GЏ��%��2�i��؛a���қ!���I�7�u��A��M����qK��K42G\nu�E����A��=��q O���L��a�i�)}����bᔘ��X�����V���F-~t]����6�r�H_�����˹F@�M X���H]X�{���\tU5���� )=�U�|��A Q�^�e��QH	RT�JD0`�1��.�����w��x��c�*�|�,�C'=�.��Jr��[	�!�^u��ShO�a�i���v�b���\T y��q���١d���0P[ 滊�l��95E)\������͖�����T�n�wW�[��T����9��3�wWƠ�4�!�5/���||^W[�d!HM뾼ZN�e���&9�\`��wv��2ӛ	� t\���L���bX�q$��-��C�CF�Qb�,o�!bC_xl$�z�{1�+p������]��`��XqwYɃ7'Xlf'HQ2k��KI�B�gx�y�2�c	����Y6����"�9��}��w��n���������;Y�{!!Z[y����m�=/K�P���f�U=�4�?>z��Ǯ׋M��oY���?� '�n�BH} �	|�ۣ�'$�����x�X��M���WH�S��`��_/���rwqӷ��-��a%A����p�s$��i3|���`�^�o62uOQ���^��/�`#�}�4�֛�վwyۼÇ��Ƃc�
�J)�°���\�s�Ǵώ�ܻU�߮s�|���"IS(�J,`�(�IW>1�|�
a��'�?��~#O���߬6�1�̔�D�	
���o���͛S�%;=A�?H��[
;׵0ڔ$<X/�x��*	�����C�@�Q4�"���0��3#fQ"��9$�O����QR���ĺ�DQg���ܱ3�c�ּ�4{�6�}�H�w��e��e$ ��}����
�F�Ĥ*������X�)Ȇ>t{u�=�\����7FE"�`��U����b�,�w���ã�h}�?���v���θ@*n8��VwV�6�Nسs���c����G���ز]yS�9 L����������	����E�~h���W��'���щ��3#��W}�[�����Ww^'�'���x{�4>�6�wW2?A2�M%m� |��sgn�4�aPb@PTd]�sƁf<��V�8Ÿ�n����
s9&R �Cf'�����n���K�N�?_9i����_��\���V����.1X-�Æ���N����>��	�(���|�}X4&P=��a�����ߎ�'��<���_r��D)$����8�1tbqЛ`���a�6̙�t����W�5 	�Ǐ�ۡ�x&��\0��hh��
{Xϼ����}5��=K;Ǆ��Wm��G�N�Y��>��8�+KR��%f�/�O����
��)?��f�|~w*��۫�g1�����a��&蔤�%}]�����[#����Ҵ�w�Wu�	��A����}��P:��;u6��W���Vk�wk`[�Ar����%[���W�G���7�������a?a�0F���+�ٍ\%�zb�����Ӧ�<�"�ß�N������u<=D�?��"�+���Ĳ3�z�#�5B�z7�g��oA��;�����^/�b	r-�i���%n}[�b��o;\Lϴ�V�x���Tg��_�����k���<����֩e�ǿm?uZ����}���d��4�vi�}L#p�CTٽ�^ui,C/���/(�b�K'�|`}�M�ARR1���7b\�Zt�y���E�_MH���>��+���5k/��7c��AL�̷��Gjp�.��C����U/� �A�aOش�{"���.\�c2��D��!B]��u�uG�,_M٤<R�,��[e�W�M���oNS�w��AGU���������SYs�^O���7�|6g�L��c-I�W�1#��&�W�ٿ<ʡ]���9����Y�KO�؆YћR�A���+V��54`9�kj×.���Nb0�[̽U4����|� J��ː(���:��i�QY�a��&��KI�-�N���׬�F�y�Զ����Ü⾇�d>��jgٚ�R�!��k�Y�K|�_�1��^C>�z�d.�O'��3P��Q������7(�#���]����E�u_M�&�Q���7�4v�����.���ٕE��ގ���ϔ�J�̂���a�3b��*�I�%��=yTM|]���2����������6��F� �Y�ll�p�w4K��j�͸DT$�]�i�>�u'5�=����yk��֞�Z�ַK�tY�e��VeN 'uͶ�9#b���st�(�Sڬ<U���@;>^x����t�Aq�5�v��b�ԯ	Ƭ�|;�6�v�Wt��7m82!a�N�s��Ͱkl�74��.:���y|; �nH�i8<n�{��J���[�ܯ=[Y�p̺����k8��۵z�m˞�v2��cu�gX�ޢ�4l��^z���y��A�mr��pn6�kd��UK7/ �n#�[v��/5�'(�n|c��ܯ;�t�G,z�&�f$�9�q�zʞ��V�_s�u;���+��?p��B�C�(j}rd�+ڹE�pױ=��/����N�g��g��]�>Y��<cm+��u�;e�뗉�qo\Z컰cV4f�d�\��<�D=n3<��/}#ێ��u�le��� h۞X�.�6mv֮z:c����٪�ǰ�uŠ�kX�1`���!�T�����H�5qP�ɀz�1��x��TGC�i�կ��� �p�^r�s�=y݇z�*��B���Ù�9wmk����E���۠�.��
i�����q�׭�A���ʯbSuGJ���x�����b
�\�i�n��u��y�WT�����Uݝ���g7n�,�Q؀��<I���r7M��vw�ul��ݫ=n�AOj�.�7v繟���h���A�û[�秱�{��z�*{��9�4^��s��ޭ3�Z
���5��8����:�7orz�q�h��u�C���81�)�nɓ\n{u�H&�����J���4v6�!�.]�,m�aFzm����C�n�����z� z�2"<��Spg�.`�tn�!8�1�qګk�@l��7kk�M].4۷�x��,�d��;�w-�:�3C��GVy�l2������ű.�p�֓L�s<���]�N۞�`���^#��&H����3��S��n���8������_���bf
ij�c�H�V����YW�6�3�n�I�0��Q��U۠LI�n]d�]y�+]KM��[�b5���l����:�6t�S��V��\�+���vi�ZX�pĵ��z��5Ѽy�hr�':��X���h�/0ls�JR�a�i"�9ܣ�����O�MM�	ʡ}���͵bnX���e���r�Z7/uS8�ff��N�/��°�����nK�O���2���-V�]��k����ĝ�#Ԑ���m8B�ݛ�~��"�Ax��v��w�9��-}�ʊi��|���V/jK2���`R��-�1�9ᗏF]��p^{��{jq/N���mϵk/Rl�m��r��]�*���tk���9wd�#)�	���}�()<�=��	f�n�7.v�ۤN;�����ݲ�2�T[+7����X��=��o=n����bH�۷�\�ݫ��z���t��H��|���q�����
m�Vz��#s<�-n�x��]��mm�q��d����4s��o9��3uf"W��Um���-iId(�	j�#�&��H��Fw=��<��U��[��p�L�;]D�f!	H��U!?���?���S��ؘ?�s���HRkݯ�w���`�v�P(H�~ �0mݚC�,o��~��"�\BA� �}��`�����'�:Q�xnN��T��h^�޺��U�lRVƤ���W���w�AƮ,k���L?����p4X�&�B!^������Okc4�{�o�}m������������7��*�f����F�)#I�i]E����>�1���O��6�#;�4���)*��*btm8�|n��9H�TC���h�!_{�Q�)��E]z������d��r�Er��`{޼IL�eN���N�|t�8�28c���9+���{[�J�1���X�-�o�:���>]���y�.�NFU���	������?:F���>>{��F!��m�7��G���sG�[3���w�pA#ЯP����b(Ēed�e�L�����dۄ�-�_>CS�sH�w_nAaovk�h�GZ&�{��D>S�N!� Y��ġ�i3x�Z�%�H��j()��Z�FŊҚ0b'���ߎ�Ai�!�ȕ{�4G8�˩��k{5t`סD�y�b����M�gi�>��c�23�N�ًE����TH���� ���!V��S��!@(�wB
#Oޠ�;F�r�x}f�9�E��~6�����V�uy�0xd��qg�Ud
,����7}o{_|??{]+TC	L���э'�
�E���ۡ(�m����v�K��jf�c���	����Cs�U۪�x���j(�F��?e���e����U�+cm<��ӛ�M͍�CG.y��p�E��']��F
3���b�҂��8E>�u�8 q�Z��k9��)�c=��u���5�X��>L3C����Q�"j|���gn�� ()J/��l�8��H�Y
@9}����G���n�Xoe�*���M�#�y[�}"e���������ic��5,�.8���VH"*��!!J�@�2�*L�"�3"E2@��D�m���Q/����~�)M�m�mS����l;���`:����s�Wl�]�|G���}��'�9J*�*@��z�ո�V1rE"(�hg�յ�������[�j�����f��������xէ�pP�^���{��[x�a|=9���a�d�	�`q���1�<ʗ�-!��%3c�@����F u������tg�2�9��
���Q^��:�lz�� �I��Q�����o�g�J+s��捇�J�������`���~ﾻ�т�~�+Fy�Ƨ�tktf��a�!�wZ�[QE��F8#B���>����C��uU,����CT����q���;C�K��/sOw���xXEEQ Y�}�X >�������7qFN�v�X<N��v�s��H�o�����1_^'��C�qs�`�C6!i�眑6�N"�!@��?�0>�7F&��Oc�Y��q�����5uzG�h�$s��7,��҈�L�(�d|��\��$��ަ~��~�O�[�Ze
�����(���_
/�e�e2�b��h�,3����P��0�	�bB�r��W��4�RS ض0F()s��l�y��X�G�橳>�.�0Ӄu9]�X��B�^��X��Q���'��R�盇��wz6��#q��s�[\�[ZĆ�nֹ8�տ\o��e��j$��l��Ydh>�-�wF:��T�����4&�И��s��7�v�sl,f��[О���o��Z�#6�f��!�8�g�~h@3��M2�(��F"21���z�y}F&|V�гu�DX�V�>߳X��e��߮��G��^�Q��2��Q�Dʡ�>����e�����Z��1��㆘� k��G�d�ŉ8���M� 2;�~r#R ��N�E��dix��ɞ�������%s����
~%�{��8F7)�����"�> !��D1WUr�7���]�w\��i��|���>�kg�c�����`�W�OS�������&P?{ߎ���σ�LR4�(5ߕ
�}�����/��԰�m���CW>mnN%U��1�+���o;�d����=��Y��=��:���9��ūl�����[���-���n�����9��C��Ql�v��3rֶ���D�ҽ�tu\Wc]����N�s����n�f:u���f�\-��k�]��æ"М��u��/F�������s��9���!��#<���M}g��EA?��4�گj�ST�,HI�J�Q��s�4�-a�N�:ٱ"D���Pth��f4a�{E���4o#��	��1(�#�>���bȌ��!u�����[[��i�9oQ����SD���X����@����[p(a�$�E@Y������p"(����uX�lC�1&��XE �E����pfZᛣ�	�s,�yَ�=ΥcD)H��B�l��o^�Cz7~Ku�}�d��j|C�ƾ�ѹ>a���Oi`�#����\�FD�-5��ۼ�"xk�]��`]Q���M	��Fn�|��ݳ��J6�E"?�, CЧ���?�6�ޫo�0���uȟo��Zo���t�_xp3�g,���͍w��`��_%?ޝ���VU�0ę���un\u�S�w77.�вZ�`�C
9�L�]��N��� o8���������JeS�r��tL�t�*����%��̏���1=���ԺS�3�F��
��a�������2�I8��,�b8 ���B�C,�ۺ"�T���J�cY(�J"���*�$���-�S%qɐ>���N9*T\;wQEV��X�#��J����~��o'�\�[9鱏njҧ|V��Z�Q����;��3��gV�ؔӳ�~�=��7�{���:?��ŷINC#B�"�.�jy��0����?���|oԐ�_��p4E��F�������&(��G*PN
hA���ZEe��Y�xz&���:�fFw�T��_&��$Y/Ф,��=ږ�פ��!�c����5 ��Р	�P����lO��]��_>�bRo�����l@���Y��O��� ��������e�\�n�h����:�m	���ũ��C	��Lf �=�K�lXJBq� �#N����C�Ӈ�0��_q!���� ��r^w7BW�k<��_���I��"i��R$�$�C��q^Y��[����w���/���2��BD^��y���{��5�Ճ,�6�{�� ��Y^���s�|X�x o���n$i�j�u��pr�_h�Q�:�U��b0V��|�bq=�d�(:́ύ���W��ᥔH�yo����j����բw_~${��,��wx�I����(��&"*(ӐRp�>���ڈ�8ٱ�,��v�&�� �@Y=%B�㽺ĸ̑L2W+;���Dg���2@ܑ�T��U4?x��װD�N`�у)W),�8:MI�D�xs4��<q�_�*;��9���k�l֛m8�xp��xb�c�F�n��7����?�۰����m���w� w�*��Cc���G��L�c�ҷ��Ĵ���x	>9�����p���7�{^��^.��A����O���þEr3�F�,hi$"*��N9�N����[+����v,���=�,=�%c3О��ZhFD�Ȍ.(RB��ȾЋ�� 4d��'rZ���=?�����ڔ~"��,��>�4`��
��I��I�P }���(�;s�R��(�X"H�F|o����Y�G`>���d�����R
?��*�D�IaX�q4��$	�� ��Ωi�q̻W�)i�Y�HL�������|�;V�+����КG��C#�>����F��JQ�s�8�6=��Y����}���W�6!Z��M=;Rf\M��Y�0u1�����������[7��[v��/8��ˢ9�7I�ZABbH!!8Q_��<�vl�˼���Pθ�=�O��p�߽�VgÑ5Wn,��D#�8Y��lo<5t`��*���%�B��~���k�G$�*H�"��x���a�d�s'�&Fc\�%� ݎ|C>�F��$'������^H�]�mwokk��ztO��P?`|0��=��)3ʘ{�]`؆7�o�50��j̈a��T�c�� u)��;\�1�%h�q�#B���}�?]���dg�L��d��ؗ�UB��M�N��{u��j���29}:��{A��M�����x�\��a05�(y3ʮ��
�B0X("-����x�L����f�Q�������5��JӋ��'�b���3��q�\�<Bl-�s�n�ig�H��U��b��BX�I ��L_|��T䭏[��6YHJ(�w��N�:�\z���8KY�M���n��X�mPq��sm�ڭ�����K�N��Z֩��s�|u�c��g�&��]n[dH"�c�����[mkM������|{�u���FC�CL�0�I,�k��{O���z�V���d;K;��wI6��Yy^"�&2��9ĝu�J�;�%��˛��	��7;Oh�j�v��\��]��_�Ϸ���~�loT�V�ǘ�it�L�K�h���cN�)í�e�m'�uλy\8;[��ܼ�P�Q7}�Y9����).8"#�����c�|�fq�N��|6a�6�O~�˫��RB�b�J`�X,dT�&�������X��'�7Ҧ	��=z��t�������zϴ����BS��5^~>���=�����K#��?�E�����q$���D��a�"|3M}����(p�\Φ4e6&x����Fe��q[薁�9>�@DBp��#��)�7����|hQX7(�dX�#��?|�N���%ﾼJM�ٯY�����=��C��也�R$�Q��J��|!�H��K�a���B��hA�{ݖxVL{�\�͹^�E���y\��l�l	Q	�p�b���<O*Zy�t�\5�����;���5�����S����W�6u�/�箌��>|��w|݊��e�{n�����`�K:`� �(<	vB����K��{�;�~�3$i*��x�τ�!�b���I�u��[d�#�b�u�{��V5~O+��YJzAw�P�+����@h��pi<9���i���m�����{g^�����?�H]~J��'$(|	#���:2�bm���=7��8�t%�xHN"�,�jy��x����)�$����V]���
DA��k)�3��O�)у�q�詇w�UF	�^��	cH�`��z�P�Ǌ�gW�.	�������D�(Pb*0�^���=F���tv�/_]��=�P��"���]"��a��/��v@�]�a�B�Q]=�z�׎ɎHp��Qn�#��άڱ-�T2\� ���D��]�j2Zwx���á>�	&�,R��ˮ�]����m&*�H�J�_�saI�V�j���؀�5���@��8!�6H�(a��X�ϼ�d��s�y�M�^�	bG_6_�6!��!��� ���ﮦ�����3�~�(+7�&d�Df(4��i�{���ȡC����X<&[��/��OI;j
��(�c'�hޙ��WGƻo��Z��j4MVg�)�L��Ť�Q��Q��J��A�^6�	%��2�UU�n5���$�ta�A��1�3/��N�r:2q#�ݏ���|���TV��� ���IP=���^�U���lm-��,��|c�R������EKjۂȼ�6�w7�$G��f勆����V.R��� n}�%n��;���t����JB1��(���B���M�4��]��IuIg���m�����3tE0�!Y9�n�rg����'i���_#cF�Ύ�]�UǮ[涫	�x�~�X&��
�B�4'@�"L�����{l�ݶ���CV�}�֩t�[��cevA�YD�AE���*M�C*�G=n�A.�+V�l4��Aza��D���0e��gQة^uLĩ���j���R9�FoN=f���j�֬�aԣx�U{4�Z��l���)sΖ�{9��{���ע����q�[	�w�5�a
���U$�i�7ꁆ]Ժ(��1������)t�e8d^�4�9YǬ���e�Az����Pd{[���o�r��w_�wwQa�&��x��"(�ω��g�.�#^}r����.��b!He(�9�@�anMk����.`��26/���C�/�)ͭueԬuN�+gA+(Rfa�c�X˪�b涻�8�N�h\���}YتZ�d��}[�A�դp�F�U{+�_z��N���7u�i��z�+WU��+���q����)ނ+w��UZص��l���Z[�.�@��`%p8C�8{��L����������C^�7a��\��UV4�i0��Y�˪n�����nY��»����P��d�;�����%�=x+�3vt�ǰ�؏.��{}WaFF����޿+V1lL�݊�;��Y�hݧ�Ur�#\��w�E'p���[2��mm�(7�=�f`Ք��\�L]�=1�w=��o�l˻2�CÄ��t�Y:�t��@P�LEy4w���c�n&����,�@��/���\�tAC�s�+D-����k�^�"Ϭ�w�V,� �ą�cHW���{ۮ��U�Ї]�6����3xX���U`:9M��ۏI��l{�~���?�lO\'0�v�.�F�ͺ<V�{N�Ӻ�CGF
��
������̃E��>�B�(�@��~��Ψ�qގ'��ꊠ�Jd���7�z���΅כ�cI��>�}�������[���M�0!h��h�У�2�u)��>��/_}�kq�c�n���L]�w�#�>%��uVhfi奲�"���Ħ%N#AH@	hWz}tcIႩ^�0Ύ�Qv3=�E�K��M�ǆ�c~��"�X��ױ�ww�Z�b�I�ha���w��HUߚq�wk���+i�罯`2�C'b ���QK,�!�Y�����\�a!i��'.sq�b��P���8�B1b�s���V��z���kNm{cv
&���Y��Q���np>� �=L��)�[n_�	B9O{��m1�u�������N�_�f���M�����#	�0i�r���o��\mrm�+���h���9���v�����65>z%��g���`�se��""��a�>�d�����H.�4]�[��{u۠=��TŅ8䈙!&l���������&�޻�}E�z�6X�����H6�;���p�d�%m��U����e��v�X̼�8�L�@�Z�1�.cͳ�m48���՞���#;���2�M�$���5�>g����p�>!�%uﮌC��N��12��8+U�B�Dюױ�>���P!�����Ouk��P��c�}����!i (j��G4&����*��Ό�d�oQQdEWi{��T]�^[mSF@[N{�79�haZ�k[����L��zN�]8�}��bq�I��ڥ�%5�����$Q�Qq��i�"On����F���TtQ�(Aa�"��Ą���4h��x���r�V�_}�Cw���c�U�C���=�tj���2���]��v8��mWm�ռ�;lJv�<��� ��|�I���n��n^Ln������ݰ�Ô�A���/�ö�Nv������8/7���V��z�W�&=�e�����ޝ9b���|��m����lx�f�:�9�M�D����dڟ�7�u�-v�.t��R�T`�=w��36aE���"�h����n����v]f��Z3W*��qs'6�&b�L��8d&$&	�j�8"�KdE*0�~�u����c�!Dz���-�+�cߍ.�����4��I��?Ή���	p��.@h
'!��>V̏�n��i�}�6||�F"`/�2�'^�}tClțe��n��j9��� �!��)l�$p#�~�XΦD��~>�HZV}Ϫ�:9K	��3��=(-YD��_��y�4DG��_���h��V.N8M����s>�>fD;��_�ZC�7%�M�4}��[��9ٍ~�C�le}���d���B�Fg�����m�{���W�w���	0�w5s�1�]�N5�[@�)���2��)�m�&��g�.��A��Bf�\��n+�]m�ض�O"�t�:KX�th����v:9B����⁴���U���P4�cw�����Mj�d�b"/B�P�=TSs�6���M���v-���2do�Q���6�p��p�28Ql�QHЃ��ܔ�|>��+V�ˉU%���	
VJ�3"�$:�v�,�տ��Y[),_�^}$�p�g��vwn�`F�bKZZ�L�~~ �.�5�.�Q�>`�������#ð��;N|mm���,Y�����(�%
L��S_{���z3l�����d������nO�&�8>=�npd���Ƃ8����[A(�l\Tk�n��i��y�+�C��,պġZ��`XK3����Qz�|$��K#AV�y���������qu��pm0�]&2I�sՔ�x��&pnO9C#;�*���?F2E�"�$��\�]r�<�DCT�C�o����v���3ۛz��]qg�K�uz��n�v�]+a8�t�{;wYK�Zuz(d�D S����������6&�|G�{���;��զ�`9��n{A 2���NH�9N�3�0<��Y��H�>%c�h�&ꌥ��g�&�'/Է:&SMXC�{�� �<�O#a�~�1�l�1u�c9�Zf$xvγc6H%ao��?a��8|�Պ��P��}�E�rS.��*`̰ҴH5Q8)��5ac̴�#����q��
�A�)%[��F����Dp�pb�Z+y��/7%n]���E��2�{�}�%�@G@��}=�|>�߾
1�I	��o���>�Q�S��R�L���Q�<��>m1�(�c�����#����$��V�(u6�����LT)�\iD�$��Az�,~���N;��h�N~�!����{t`�`d�����栫CeZ*�������󜐲2�j4�#>���cϭ���ݍ��V�i��+��Bv���UԼ��/]n�F�h�����+�F�z�PHa�d��B"�o�Op"���*���᱙x_I��9�3s]��� P8}`��udL4dR@⒩�XFz��=�	}3�:���9~Kg�����:����1:��:��L�n��b0� ��i��TF������ܷ��t�l��b-��b
��QI�X=*c<|��xN&�U@������Q����s<���#nHNS��~�}��J[���i��֊nn6��(��Y�������+�}��ѳ.Q��5�^b�4[=J��U����I]~�-�+B��xo>%|n��a�*}�@�q�ޫ̊;�/�{7��f&P9�U�O��y���%����F�k �m9��0��C���M�(�rH�owo��N.5#�x�zM��pE�wn�]3�7k�aƐ�8�&	0 ��5EU�e��\�g-�&���>�J��6�"hg{�xd�Q�]l��\�f&^�Ԭ��q>�`���s����E�W�JHL"<9���>!nD�:n�C���������4$w��~2��k�c�[��bH؍�k���a�S�T��>�\�pχ�b.=��>y���xfpf��o�Z�>��������]z��8��]��
4�m
�/rN������>��*�X��^}��FX�y�}vby߫4�|�0� Z��h���ԥTb�V)���g��愳����j)6Ũ��@(����K�m��;]i��P:E��I"�`�rJ����la�+���I`��}�V�\5e�,G"�ܜI�S�vٮ>l{�ă�>9X�x�ʁ�H�q,���Ģ�+Ѷю�rɳ��ێ� ���B���u�Y's���l]e�5�V�F�p��u��0N��.����F�ݱ�Ѣ��_Y�ݸ;���F;E���p�e�ۉ��{$�o-�)�g;��[d�x����WV��i���W3t���7[�|�<uQێ:P^@��s�Fo#ɸíw;&a�tF�a�d�w�7��Z�}Cpɹ�X��5*��S9�d:&�U�E	�0X��lZ�9(m��ݎ��/cVcp���6�P�J�Z:F�H=�����[Qȑ�Db��1�bK�;�'�j�z�]���0;L��;^����G�'�*o.+w��'�_� � S���'pH�M< C�!�����-�s��!�I^ğg�\�8�G��[��9��I��o�]����]�s��}}��&�s-	���R�g��j���LbK�r��`�ۡ;���ą��=��8��$��ܦ��Q��f��jγ���P̰��t�6!�[�gIxs�њ���IP����]�
�b�q��*�3��@�_R�lw�qI`�4}��xz�Q�>'KvZX��q_�������(�s~��,y���3^ţ�j��m]�f��ֳ�G��r����[ti��n�V��=Y�Ӻ�)��H�	�Ӂ�Ѡ�O� I���՝a�.���@�c�e���U}͟g���l�B���Kiȕ���"��6L�J�H~�vi!��~����x;�V�)~���'�8���7�ݣN�Z���طv�8~�?/
]���hv3�o���:$��x8ˮ�٭i���=��AP�A����D�NA#nK��~D�~��FeNo~L>�k����C��ک���Ȟ���#ߡ�ފG#p(�eq�a��w��z^���dAGf+O�ٱ��}��3⥦�û����cŎ� FvZBi����.%�҆8�n�׮�4���P J"��A@Thƌj�����I�PB@��c�]��������40W��>CCba�3��fm�ݽ������?��H�^֠�j��O�L]:6��g��s��ӨM0Q`$�%��J�|r�5����7w1��Yl��!��4!�|�O0�(���"Y�- ��J�D~w�^��M������A��x�i����
�Ӎ<Fy����31~�����Hu�4;�ݻ���l�x�+�L6��WK�2DE�bşIsX5��w4��<��u���b(�#B|E���~�Z��8x&�2���c�(��SR�$���33��3a$�b�9C
�"J�RH��$��1S���'�{c�}���U�f�3U�ځ>ƴ4E�	H~���K�tp��	��q�6���I�$a���hP�<A���x}	X-h�o(�(���"}��<L(C���x:}(�du\�>^Y�a�"����"��7蚈�B��� w�K����1�[1���%��)"�H���;�'�E\��Pɪ�~��y��e��#2�L��?����y�{C/l�u�/)�<Q��:���i�����]��.Ju�����߯����a�$�764 ��HY��I	�������>�
@f�"w�����P-)=��Բ8!� ,j:�#	H�r���>C�{]�9�ki��Xc��s,��&���6�)`(E��d�b�43�ȗ�/�*��PY��{|�F��||��8|:O�	�~r���4(0L���H֭{����ݼ'c�w�x�jO�q��]}wV�JD�p��{�>�xI�C	vɢ<,�����`��Fv��K��ߔz��J A�>�)�DD����"L�1d����+�����B�H�d���������g�>wxv.�*<��W�5xK��j�Y��6_~�M��-9���	۷6��u��S�}<�#�8�*:2W�(@��>l��ݚ�X�d"�1W~�V�Z��CU�U��3��Y�}x���YR���?�u>�����K3��M�mi�U�ٮnW�T��PB3q&a�y�e��m��2��\q��� {:�C��5p�Q�gk�4��o0�f�'q����h�Ͻ>��,��n�r7�,��{�l���ǹ��e蔸���M��(*@>��c��1����{۹�Ck�+��G
��6̎(�Aěw�3��;��g�(pH��Ϙ�ֱ��C7��bm��T)� ���Sįa������a�fH�������`�s���k�]�b'K��F ��E�2�$QA��w;��}�z���`M2w
ޡ>�B[A1����
�xI ��)�03�}˼�s�:guf�a��yt�C����9|;To'��YCN�X�/��sw�c7�j�3��dTP���0�^L*!�;-=8�SvC*���f]�ٸ��D�^_�ժ�r���6��鶬�%fʱG-q�(#צƙ��� �H�W}�g,��"n�����3U��ik�>-].!	�R�[N��Y�LH�k3�b�TJ
B!i�Tr<(Gh�t��@�wv�����~b�0�0������v�b��T�[�](����rx�lY��5�r�}���j��/͵���,�U�T�m�����&��Ym5�u6?D����.�(����wӛ;z�n)�n}-�6�U���X�ֱ��-���ӞeXQ<A_ɚ?f�+�E�7�L��%	L�]��s����OqK1ќ���a�vA�L�^�h���_t�ɘ��s���_r;��/ڴRՖ���D�qǅO|��o�;/�>����>]9Ӳ^P�W�ܳ��ؑ�b�YO�����!��r��>!�r2�5A��2Ȫ!�j���H�3>Cr��]��9�2�Q\ɷr��\yY)�N�t�UAX�Ck��W��j�.����Y�֪���թ���Lf����5^���3�!�(�^5SH��.~Hm�!>��z����[�a���m<�b����hZ�*����I�T�� #�8}�,� ��a�K����������{�m���\T��ϸ# �@||���O�|*�� ϟ���h�B�٣"��(�(:gf�R��.���Pp�:,s�ύ�!<f"!b)	,l��cp�;[u[5��H팍�m�g���$J{ew�M*^[A�孕��ٸ�>�⣭�1��P]�v�g0�*byESwi�>msv���pL�Jx`��n;M�PY�8w�98.F�O��ۃ=�գ�L�bl�B�{s�tY��s�_)ː#�-���2g{k'���ۃ���zPvm�5�dG�!n$t0\[ �}L��x��k�9\��vQ�z;l񣓔�8G��qE�0�.��\m�uv�z���s�W��\PF9R�n�{yܙZ�b�[�g�{$x♎v�W��x��Ʈ���-3��:�ݞ��f�.`���[�y4�n���M��:GEK��8\��i�s�
&��+<M{v`<5�;��2��v�8�E�gE+��볶6��qr��2^��|b<�ݣ�b���B��m�\������qqܻ�"�n�=c�+��f�������[�������G]�S�Jι'/Hq��^T��r�S�W�Ԕl�;fyɌ;��Kv5�8��.-�C�n��KŜ��{qɇ �\�n�t�G=�pm����7�xbU�{u�O�{u�d�q�٫��7m������6�I��V�ގ9+;s>����\��u�.l۱k���n�1Ƚ���0qí��tO{+��x���8;Y�qi�a���P
�(r]�[�<o!�u�.�ݶ�s1��+h9�8�GY�W<w2fճ�q�F[���b��U�;v�M�M)��1�=����8VA^ѣ��)�r�e����v�u�������
�Ζ3Ӯ1�Z"'�M�\�ι��>T�2�ݺ�j�.���&-�ݕ;��]������������b�v�b�6�q�yy�/I���j��9v��8��j��G&3��мE�Qy�Wm;Vv)a����Ռ^��r��	��[�����q���x-�;k��u�tF�ޓ-��4z�.v����Z�\���U�;7�	�'CT]��ܼ[Q��c�Ƿ'O(��G�����e~�������I˾*�/+�,��//8Q�lJ�.�n�M��ݓ�k�L�n�v�7K:��8�^Vr���[�7MD���5q�a5��3ד�S�`�Lg��OL��-*���moj��mP���k]������T�%_�ز�����mj�U%��[; ��c��s�d�W6�(^��oa����D�{�&,�Qwg��Y5�8����/�%�X:b��]t��!�+��ە��{!�k5�f>�"-���Ǖ���_L��$��k&]�vjW3��J�X��Pk:�_o����ݺ�.H�]�	;�0� q��s�K�ˮ�����⎸�db���5UG쭽�;b�2&w^8x��G]��ä_W[m�秓�W�����cn�Jln+S����˝��gn�{cLeknYvvy�s\� ��rf\�i\�v�c�j�t������8+;k���-ݩ�2�tƆ�U�Kz3�/��޶�'�������h���^����>}ʖ�+k�KUrQ	Q̻�$�����u�U�O�lp�d��<p�\;�����,E5�D����DR3�H�-��R������D��:ˢ����gk�\.�6Kg��.v6�W_6oU]���|4����������3�F�Eƣ��F�P|}�@�:�_�}��BΟ@A�cwx�-#�J(X���M`��-�L3�����Q�a��M�[����~�B2H�e�B�DO^!�{e���7>g�4���فs/��oa�{Ƭ���,/�q�}���e�7��\&IP�#u*�B O;v�d;�:��8�O���!L����'GǮD��f��2j!b#"�bb��桮�Cj	�\@P"�;6Hdح}����11����O�=^��L��49�9��n���a4�H��i[<%�3זy-����Ywt�ی�j�-:��\��2�Zl���s��R�rl�r��~~�o�??7\[�]�Rv�k W��{>�љ���$�;��)2n�"[�w��wד"
}[�f�W�?1n}}��w/�����E�:�~Jgo�4���*��>������`"�5L�.	 ��9`��J�M�.3��*��H�P�",��\󭜤ba�;���	�ݝE�UM���Q���Oyv��w�w]s�p�y���E�,��(F$1s��R��r2s	dP,Ngd����W����r�S�R8�S����0�>���,Y������58K�1K�w���}	 ���5�@_�_��<5��q����������g%u��O�μj��
u�����4�M�;���y�m�(Q�(��bǴP�o���|����Tt"i��|�Wx�W�]�bVM����er�받M�1�����=ʣ&�/ϯBĚC19�z�;���~��o��7M���,�O�s�s#]�yz�=]�������A�1�n�Sۙnmq�IQ��=x�>����<G�D��Cc0��I�i$�r��û^f���N3�xn�`g�����Ӌ\7�Rb�e[����i��rNُ�e(�s�@�a�~m ��'�8I7�z��|G���{<L���g�[M�$RF�p�C���
�H��U���BZ:�\��d��H�&��)̒��Y�t[6�Q\A�ՊV���2J)%\��~'O�#�p�0��i�hf�uAH}�Mֹ�b����v��.�&�`����|,�6�6�Q�P9E�[��L�|fr�=�)sB[40X�����m��}tbm�N�0�U"]i��9�D#CM&0�$��KI>)�<v�דVsY����2=�}�0�cH�	�E(x�!�l���}_�(��l�TĿ��m�e'GL7z]& ����1����q��UWص�A�.MR�ɶ��� î�rz���:��k��j�褛�D�?^Y�$�1��猪W2�fG��[: a;�6pe}\�\���X�θ�ڽ�(m���1n�P�\ω/�dA��q��m���?�M2%_���u$�Y1��ʓ���
/ׄa
/^��3>+Iq��U�0������wFM�:0B��n�%�q�"R��0������& �����q[�督�8��̦pN	]{�хN'�7=�}M7�֩�BcQ�^���~�����$U�@{{��3>Ht�@�!�<>��s��u�Og��|Z�I�rEVZps�F9��Ϟ�=�ο7��[_����Ӿ̲4��A��t��K���C��|*/l�9;m����1Ӧ*������_��kth�ca�>V�X��Xpm40�(���������J�j6���9!�(a0�����A��x��)�"$�$�M�f �p��v���RFmHrGq�i�J>L�x��}Y%P�y�}x���>�yÌM��8&���O�!���������꽎�y��������x��q�pd�՘a�q���I��!�����q��/bm߾�	E����c\T3(W����S�f���9�Jy����q��ؾ��De��|D����
G��O��]�wF-�Ud��G�w�ۛJ�t`�P�n�l��'R�Z������pOgeu��uW�*6�j#Y��'znkx�c,d5���&/qܻq��O�m���w��;�7��V��o�FC�4���� ���R�u�{_]�dF��٨��I���'ͰLQ_�(?�y���.�@�hʊ��R���$���;^B�^qfJI_��rgawݫ�ސ�Q6�~ �^�m�
<V;C͞:�h��3��������y۩��:������j�Y8�f��*��<3�3���V�nM5��8ᬍ8��m)���&�h2g�7g�Z��[��>Ty����;p��h9�͌�m�ąػm���훭�����jp�n;�Κj�l-2Gj:��9�$۴�L��]��Ω�l���I���ƴ�DY����w�I�<&N:'`�C���j�����H��AV��D�i��$�mޒxqZ87i�]��s���{	ѵ�!��1 ��KEÍ�i���F��F1��0�e���5t�O&��ͦ��O_������m�X��_�
E����|�0�M��ɜ�𖞉9Bv�5��rl/��ى�!T��j�u�l�w��H�03�9���R1�E��u�"��{|�`����S��1�l��
��a�'��a�e螛�`��a��G��z���������m�ɉ)�HF�,XD^��񲌊{����h�5���-��Wۻ�;G�� i|u$&�n#'�0}�<��|�lȉl5q(�xz��o��'G)���.�ݘf��J��iwF&R,���K!��45���p��r@��0Q�Wnmm���J^�=�A�m��3�eB����J�Nn��fD�O�v�-\<�O�h�{Bt�(sG/ͳf�g1]��b��|@��,��A�*LY����Ɂ�������l���4���8X=�����������0�R��!�@���:��M��k�)�A��<o�Sb}4�P���Ӱ$��,A�˚������ ���4���T|!r��9�0�4Ƃ��I���X��A��Km�Iy�E��`X�z͗X��u�G�/�PY��ߚ�>�|����I#T�Y�у{*�)H ��)v���ѭ	$������`���>��Ϳ�#�v?U0���zʨQ7&H~�in��Ąl1PIHg��t����|�����+F(������=fzVx2��}D�V�B���$����A�d0�@s՜����P���/5�L���D$�Ny����Y�kI��$�.EH~��� �o��P!�v�u�Uw���'b�@�)������{z�1g��w��EFcȒm�K"�>\�����W��@�:��a���-[86�ލ��Y<j(����(gO���Ă9 2)LS����������}�������~�(��of-�ĪX����^�X��ު�[����E4a
Y[ NI������Z�`zH����" ���TH�VO���w^���������cw8�GZ1{;b��ģ�~�>�K� }�)!?PN(؊(�j�#A}9|����x0�����i��go�yn~np5��x}����窽u�s�9�tպ�]��(�.��9���v��\'=h����b~n&�3-�_��|-	�!iD�G4 �G�Ă�(,T>����9��ɄɃ�$ϼ}7D��ۄ4Q�ľ�������>��$#A��F�|���k��ƃ�94P�3���<�nE�$�$m���B=,��l�p��}���>��]�r]m(Ǹ8�J�eDdHR"Lq�\��\ >Z���ʍ4T��E'���{�MƱb�l��h�""(�o��F�3�s��v�멁O�?e���<�����R?̍J#�9��N\G.c�N���*�%Kb%
dL�T�)$AD0�K����zIG� I! �A;߯���/��vak�",!K��&���˕�26c�Vnu��_�f�9��Ɔ���@����ig7{ȋwщ��{u��w�Ӄ=klڿ6��v����<��]S�>+z+���M���躃kM�=Vwj1��ܼd
�����Ѱ�&�\����B���~&�(�/e�4������˭:9���
E��0�<�������o�C/o�JQpkaf��Ԉ�ٌ�
I��(}g�k��kjh��i�8f�Q�٪���Ń!B�n�����#֩|5�Bn8�F`M�Tr±��&P�<�F��1���[��n�;neۧ���ga� tdY$U3�_`qt�-^��lveDFIF�.�u9��{��Ӏ����{��L�`�qۥP�6Ea�n��h�O8���?~1��;��pq>�q��su�Y{R_���������BĄ	$����� �Ѹ}!"�Wu����W�t�wI�MoT">$&/4ř���V��"�!=�l�C�e{Mufbx8G��W�]mv���#�kZ8ua:i��ƧK���8��W1Kv]vP�[<LK�ӷ\F��}�m�����V�y������wY�쎯:�G<�v�f�%6W,p�6�]��.)��^�S�HU�<6��9	��/�aۡ��3����3�����q͠���xκ����Du�1Q�,�� Y�C��9]v�R1�q���wUړ�^Z]K���9'I�����Bs���nH���'k�Y{c��e�v�<Q��&�%E��&�u����HHȒs���Ą����#��g�I�`��������]}��W��(��*Zi�{���
�I?oy�a�F�tS9�BoԸγ��\�o��2j�Sـ��~ ���p�I�����2�r�\j�=���_�ߵӣz����>���RiH�HjR"�Ab��A���=��x<9T>:K�)d>�`�^:�_XBGa��tj�,����=;᫬q<;G�}�}F�C�|��g>9UU��������?'���p�����V�H#�B/��Y_P�j���A~ �����?v�p|2��'>0>���K^�� nL��+n��[jn��u!�7���ĸ88��1&��$�������1��I�X��\�`���"��C�����.�f(���U�~3�`_}�i6�n;�B���W�6����'��}�NJ��-�:���Ty�AÎi�O8(M���?{߼�?F����Ŀ߾qR�ǿ7V��>��E8Z��dd������\�5�}�|���ߗ��zcb �-$�#/�������8Hb!9��:¬0?��~%¤n#�6p��4�P ��u1�V��
4õ畉Be�{��v��C�D"
n���	��������+�K�w�e��s�CF7���ѭ<]&�?����~H���?!C>��� �c��bkk�<��r���rR�M���wY�c���e%xz:�G_��/#lHm�S�K�`��4�Q�x&��g���9��b�E�Ǵv������E��߾p�!�@���Tn�
K�:ఏޠ�w�5��W�Wk_vj�����E��hG����jC��,T���ݤ�
�k��#����"O�R���5����3d�ִZ=���"�@��ᬱ0�#�c�ɔ��U��f�d܆GN]iGf(�e��q�]U�@�S�U]ܩ0�eS�Y�&����"nUf՝k�^{L�!�.�֔aǮN�����)>v�0ʆ����j�BN�k�'7h؁�Tf�:Dtp��ځ��ƉZ�4�0~�[�0+o̜��"V�f��d�qS�,��dX(��.�פ�Q�Eg��f�C�̓��i	�1n }Iw#|�%��%Ǝ%X�s��(b�u��$����9��X�Su>���NZl7�A8Q�>,r�BrV<U�a�oM�!��񡇏DB3���x�2�p[_j';8�$9��э��Mk�)�U5�����(b��4 Pr^9H0�t�6�=5��I�v0~�dOQfƴ�
����A�����I��)S�DF��f�T|2+4�'�Í�U�S5_P��.X2*d���X����]לA�'f]�1V�4�
ۻ�/)1Bʿ4�ׯ)Z4U�J�$V��FдU;1�H�
���6#�5oeeYa$x�
�Խ�0�k�\�E1�&�3��i�q^�-�R�Ua��9�bWh���T�L9e�;�ʤ3�%��XJ��K��Q@�T��B!J��<r踵�~�
���l">�;��c��]�0��W��7轸��ig��rNWŻ����[��b�Y~�!4�,[$� I��H%K� �Hu+*�2g�v�Qq5���.Y��V�-�)�7nI�|��G���Y/�I�C�r�mf�:��Z��݇\�K �]n����o{m���]�n`Ȏ���{��gE|;2�mr�v��$M�y��s�x0<�νT!�B�XG<�_��v�m쩬+�	
Pu���m�w(�w,��H�	���/�)7J_�k�ة0���ٕr�R=�W�l�gUE&U_+��6���r��tʛ�¯�Yc*��`�:6��z��!��'9K��Lov����*��Tt�3�U�3z�|^4ݡO-����٠��[֞CF]A���C��<_! &�������=�A�H�m��p�t���_�c��V����*h1�[b���	ߢF��6��A��k��F!�M�Yv�o��Q>������yY�ٱ�":>��V���=�&����E/��9���o����Jq;v6�x�v�ͭ���Kٍv�*��>^���u�j��EI����t�����3"&�!q��x�AJ{���rϣ����y��o���RB�w�-?`���*�l۝譈|=��|�q��g�	�D\X���^φȿ H����o�����R9� Q�F�q!w��N.��	�'=�`��+�@��빠���$X��愡��Kk���pd�>a3��mo6����F�	����s���X�-�}��p��j�;&qES,-��	Z���f��꼱+Fܟ��+ͧʳ�T����qiٽ�NZ���_
��Ҿn����1�d
(�xjEwr_�/�,�~=R����o�Y�E�o��"�l�Bɉ��ݸ�0��߬�gi/�x[�W^�\I��k����u�L�c1@��a�I/��;̐9&�bS)8"^A�~����G���ꯎ`[_t��� ��~�m�Fn�[�6��i�n�o�3�A��G���hVݟ��j�� �D��kJ�|z��@�~���²�?E@_�u�H6�)7R���� ]��@���|��n�o�b\�D@T�!��"d���{����Cf�7�1��A)3�{:t6܉�	jK1O��ڦ��k�O�ouEo4}>dY�����嵋N�~������=�d����J��0�*��.��x? >_���V\�t@ա��oQ�-��wy��}.ϯ?<�����q9�^���(��V�����|��k$hX�-wN�Dp[E�>G;�j���M�ґ��1db����y�ڔ�u�����.ہ�Iش^%���\g�K��P�n2�j�S���{n8��Z�a�� a�Aq�Fkn�e��{3��V���a���z�U�֐�poH��]�bn�����m��l�<K�ۨϮ��w#�y�;�vx��v9��nd�u��N�&�]����x�F힤0	��7\������M��Sd��{3iW����]�����כ��#h���0R��[tfƞ��]�n+��:�A������*\�uS]SXK&�.^>�r/X�{�3��8s���FA�|���L����y�9�>����|~�R�q���H�P>g����4��wf���@��9�I�n�Q{�4ZQDb�/<�=���f�F�E��j3(�I`{�G���`������Fb��>�>���@�������4�O�%����%H�i���B(�U*5b����<΅;�}w�&P�>!_sU��I�7cc��~��,����% �|>�{���S2�Q�uF�pѡ߸(K��V/�/xoes����������|����X�^�O�T�0|�p��ci�MU�G$y�[�89��\��۳��J�G��/�S1�jG���#�Q�����1b�����x�7��cx��7S��c�f���A�_u�����;{���t�3�����������#&��"��1��B�i��D�FW*Ɇ��Ō�mD���TW�������Hk-Uw+-�4s��P�z_$�V��q^�D�m�EV�b�O���3���^�u˽׫B��h�c�g���Qa�]Y�-V�H�C�'�g�|���,}��k:Q7�8�Vf����Y<Vwv�f�B��!�bO8�P�2���e�/�J��X��9���;�divX2`������+;���p�[��"m��h_�_rQ�������x���2�>��A��_�]��x��o�u�ʔ��o,3�F�W붬<�=��I%$�F���\<y�|�e�Z�$$ɱA������m�i��U���N{�ⷬ�}��o�1���߄�_��]Ew����P��k�O�.�mt���x/t����+=����>{�����^���%���������;�U�y�okc����O���ߥ>d9�A�*u���/4dI��M�<|��I�}�n�nS$"��?\�P[|��tuR��t�k��W���e#K_�Oz3�i�èE��bX-��=�_��=~��r���<��u�������c��U�#��EP��!�ř��羮x潿[ϛI�h43Q1T"w�}���w�j�=k}V��4�w�
\��W>^�\�a.�5���co`[n��Y+5�vgt��-��r�JY��✴#%���O��,���P�[������#������9ڣ]b͇�xǜVu�.�h��A��9^��?��YO蔐1�&�i|.���~�]]�\�%��bF&�����P��'`|Ϲe`'kF��co<�A�eFAAH��E	��묹�6~���c�/���Z)8�V\$=�p��Ԧ�X�/~ =+�w����H9�Z�݊��mF\(6�nrc9��� �>�F����h�Sb&�V�\q[ٛ�:�E����4��#1+/�D�JEk K��u"��A�ȫ1���u���~�caOs�f��Z�6�#��kr�xX�^��X��ĉ�U�*�9o�)�>����P>�;��b�����%��Bu.����2�����~���k��ӳ�WWtR�?��{�9!7J5iIH�\ߤ��K�\�!M��h1s������
`�)"Y��5�˧:�YwRϱ�YW���\5!�`�vr?�.BdH[%j�{���q�~����x1J�]}�� ޗ߂nQB
o=��㾪��H`ڢ

��������gY�n�I�,8C����׈�=a�w�H>	\\�"x}�ԍ�������ߕ�����O������s�)!;��σ���'F�hw�H����Lvi��	���睦 0�'�MND�6C��B�Q����y��A>}�T���~�n����%%Y���z���_ϛ���wj����,����R���SQE���ϝƫA�m�������֒С��j�%"���9|`���u�� �m�z�r'jg�� �n�E��9��\�]�C.u�k���;n��9^՞1�;%6�y�]k٣�AW{�;c��];f����ǥ��n��<�k����c-�v�цd�grdC�c��vyS�{��Yg��x��:�<n����Z�N��F.A�@�k�`����<��b�;Su�8�iu���P�Λv��Nje?��<�����u��Lӻ��L�J�I?;pv��6���KZ��=�n�ҧl��<�nղ֭nw#=� ���w�ߚIr��ءQ�|9hE�ޥ����W�_#^���o�V�Ñ���G��^���,��cH0Ԇ��T���|�M�'ē�0D�RR�C4�`�(�������ߑ'����>:~?�rfj�!�E~��퉄��X�m�\$hy��n]J��N(F�,A{��ϱ��fM�G���zۑ�sX��p@1�h�v�r��?���;�5lOG)H_�m�"���P�>� �<yPZ�Gq�@3�:�JKJN"��@"k��#nG$���� >!�Hl钎�f����mO�5�tۼ�<]��sU�L�����S�N��-�m�V�[g�7a��::,���Zݸ�$��i����{<�I��|az���>+�u��{���4�]� �R{�6*��iVB��~l}�P5�����M�8���~h �1��$���)d��""(XI"	(��W������/.�yI��<m]�gy�P����[����u��7���Z��5˚جQ?Zx}_�,}�T?o�`���D�jT;��c""�FH��a�������h��W����/qʬs�kh1Ub���QY����s�wr��fj�}�;HL��2a����lZ^�N1���h΢{et�Z�M�]`Gx0(�Ué��I�#1��P�C��z���5�h���.8K���>'���<�)�k�i)�H�e�r#=�4�Nz��B��؄Uݛ�s�N]([��s���ߞ���Ӥ]t鳿1���q��?~�~K�Q��2N"�
H|��P%+x��-r���������A$A�#d�UAHW��$K�>'� #f��2�����<˥$b#>���G����<n�A��ߺ=���Ñ>����}/���p��iPg��߿7<|Q{�(#�
���?�(,I�0�q�PHh�PI!��U܍A�C~��u��Z]}.��9�Y׭�΂pVn]ۑu֖n|?��?�5�(�Ӿ+�$����L	*zJuA��{�+5Y�yy~�)��F��. ���`٬��#7�{���TV�w<�.�M%}�z�_z�fܫ�-��+>'z��_���3�~��w��Yi��e�B�������p;�����/k���^�ͧ3w���@�}<qé��R�:�g;�������f�h7��"C����
.~Wel�U���_�����ΟOQ��i�gW'l��-$�0eT4�Q�~�`\�㿜�|�F�h�Up�F�
�PE0�3�x3P�hnX��$#]���Ua���'�l_FˆF!nJt�$'�'k��XӯS;��y'�����}>ɿ)PL�c�_)�A§dIp'$MQ{��"WZ�*�ٖ�� ���Y�|�}w�
�f$��^����������������D%A3�3��Y��y������^�%�������'J���U�a/j݊���[��ԙ���6����xO��r �F:�J������.�x�z��|�@x����RWj>�>�� G�$@>~ ண�pF#�:�*c��%��ݫ+{[4�U�\=t�����n�������~����B(c,�$�6s��u��4 R�Z�C� ��7�s�]�a"	�~j���Z7x�ڂ7�������z�*q�����(��ޗ��`���4�I�
�$Y��b�#�cV'_d����$?:�_`�zƯ����H4ۍ%%@�����|J�>�� N繡/�wFL�?ae�JTW�w�^_{�\_�~`�Цˊ@�qD��}�|���l��־���~&��� ���\s==U��b���������� r&��4�_��{�o�n�5�ϧ>��7SN�����P~��x)ǌWA�����O����ʢ�.��Yv���Y=.�c�������'��v]|]�d���������RC,����jE!j�3S��l����(;�ޜ
�$ӻ��{�;�
�.Hŷ����Ӏ��ڟ%�)K{�p��n?�Y��
ƻ(ɰ����������"B��qJ	��������k�&���t��_��}6��Ka5�HZ���Rb�f$��+�����xřz褫�06D|��ْ+��h�Zojf˩j��w�"Pո)d	@�y}�2�؆����n#p2���>��UUjTk`�	�����©a�a�R�3w�0��un��������*�&+-��v$	�幸�ɕ0��}J�A՘4��-�{m�K�2��0��sQ�e���4�\�
��Y�k�:���v���3����~xªl|�!,YR�iLl���"ڣ�M�!�O��-V��K�R��O�mܲ>�s���#1�S��}ٓ�>�+Ԫ7���)m��	�D���M,l�J@T�+��,��^\MR��̫�Y���<�n�/�[�+I�	�|�^]Z�e]-��#,�C��NUCz���8�v��d1�/��ղuc_-M�"��� ��c��5t�Ws�3C����{�I�֐�{���x;��� ~�∯�@$���w >�q�o:f+��bgs�U*?)�-7x�l��~2g�W�I�IM�d�<8.N/�_��@�p#���d[D�MB�IO�@�1�(^jE��#R��U޼�B�ԎM�J6M���y�u��R:8�ݐ�μj�vS�f��R�wnt"��U���zn����ccz^+�vz���0iڑn����ܯp��N�m�Y�,r+�9���<jmRl�2�zK�۵��p��Ԍ1%`^�N7��8�]�=IͲ��8��ͭ�u�x{F+u����,a�.p�n�3s��L�k�u���\"<;���f��<���v	6|��v��y��6v��-�yWo�n��N�x-^��i�v��-�Q��ܨ�jJǗ�Y�-ms��j�ttn�gǔǁ�s�'e�4���4
�Zs9�\;kn,p
�=�Q�i�=o�����n�;3�#��#��zL;��t��Jr���aG�8Πɪq���<�#[]�t�{[�yNt�lF��X��t���'z��źM�N6ol��rv7*r�������hɎW=^ �7�Wr��m��:4�]�:<�kUm�!CY��9P���K����7E�Lb0�0v�'��������	�`��7'7�Q��k��4�郎@���-�v�z�<k�Y��k�c�}p�#�u�a��v��a����+˦N���2���068z��7=���k]�76%5��N��f==&�m�g!�*�l��S��;����\�.�����;:'�5��y�ݣX���i�(�kz��t3e���e�/lsMe��\�ݎ�����c[tyvףro>^ܛ�t��k�0U�j:�qk3���AW�7�{��ۙ��]�n��W�M��-�A��!J�� u����S��� �7�9B��.�4c��ϣv�R�����{�p�x�4�m�zN7v�#t��U�{H�:��g���疘۝�A郃^S��klvy�/W^\u�����w-ό��=nIݯOe����h������ٻj��EtxO.�%�kݳ�`;zgs�v���Ż.V�9��#�uQ7��-�0u6�P�3�t�2=��H5��<Ώafم�Y�T���y	�0�r�*�5����fgd�4[u�En�#r�ϲe�VY:���Fn��:�m�f	ْZ�^��y�5�5�d����o��3qI�9�k�j���37z�:U���ف��Z�w%�Ϲ��T޲��ٮB�v��31�k�mp�����4*��n�h��/��� u�ͳ��tQ3V>��f]�nQp*+���hbW�d0�e��B͍��{v���ή�ԭS��P�u��.�/�f	��94U�{��n���A�Wyq�a��՛e!��f��<��hi��k�C7C뗤���ձt+�g�m�c�]t p,��A�����疹��-��rK��n�]mt��֛�R�FE�&��)��]��l���w:GMŔ7����%��띋���Ǌ��ٸ�{\�˫�;�������rکa�^ݹ��1$��0�En��X�#m���nK=��vS�m�j�"�cn2�u���ˆ��&�7C��L~E�f���D�:7V�ݲ�e�m�'Uw�VTr" �h�J��=��nv����[U�M�b�n�mN�	[_s���wbF�.H�"H�F�s�}��G"}��Ϟ�ś�Z�Z�+�}\)��޺����F��ܹ,j�m�_��bH�a��`�DSD}�������^��7W��Ҽ���S3��ݺ�>o�^�����:����i���IT�����<���~j���Z�J/�P�7?N�id��&�Ea�{��i�A?�~�-Hd����0N��Γzl���[q�����U`��u�������^z��K�l�(���z�O�ӻ��`���4��d�	4���11���^E'H�泛���r�w��>��5���1>{�?�q���'=v"��[��)=��qͼ�]����=K�4(s�FTE42�G;I�5m`&C�8"[ف��6~F~���]�T���ۛ��D`VF

�_�2^k�p�ۺ��M��)�>� G���!p��r8�r(�G���bϷ˽拿m��"���)~��A�l��r�d�-F�m�����y���{t�Uu������UT��J9z꫕B��̣�vd��cO^�9f��`C7W1=��%�;�z��F(C�>18y(���)F�rBYx�1��tcg������O_�cቃ���=A�l����x�x /�_K:��Z�3R'pHm
���ݏ�,R�K���� n�:}�Dh��~���d���/�i�3������/�Mʐ7%,����|��B��EN�x�T�2���B(H�G����[���G&:]X���N��Q���s���D�/����8�V\>�Jμ�q\�q&�?�!���I��F��x���F|1gkܪ�fk[眚�X��@YQ�5}�pmOD�"�R0������Vh�]q��^/G"�����X�a���ɲ(o`U3�
�����G�c�ⱏ��&��S%澫�=�e|�D��q�#����+೪(~^lu�h`�.�A UpY��A6e��FC�8�-�MUK"�2L�����E8�3T&����-�G�Nf�y�������"�gL;��E\�o����kj΃��OB+���ܚ`���h)T��v������Ѣ��>�'��B��Rb�<s��_����D�B!���[c��ah��ø~/0&X��\����l;x�Q'=��o�Ϯ}��������^`���Լ�c;�'�e��7ߚ�We]�R�K,/0U�NyL���)Sν2M��W<GF�l��:�m�տK��E�`�#RuQq�����_�m��^7��l�������" �b1b1I��9�7D���CE��f������ς�Hp�������M�[r�$׉'T}�K�|>tw�����A��.��#��:������O�߇<X�{	,��.
uQ_�Yc��\(P>2/���{�j����\t��fph�~�}Sn����;�����������ᴖ^����!�_\��������=�{�}�>�wu����j����>��8.^�lyug��^N���r�H)e����Q��*)!�ڬ��Y�n�Y]{�O�+�"�����˧���A�cֆ��6л'�{��>�/��8��R�⌸$�,���ak���)�Vp���z��Zs��j,��@��Hp��#B����3��(#���RfmM�uW�J{ûbȢSDTX��wx��9~68/�_��'����f
*!���N�� ׻��G��B��)�"7�x�|�G���U�#=<^�K��ֺ�'�_�z���:7�Dg��|˘�^V�[ݝ�������QD�z���X�����ʽ�&�2�s�(e}X&}�0|f%ahvw������ߒ�@����|�_�;%�pq�8�b�H��9-����{�c�}F�����}va�u/8I_�F���DP����f�~�Ч�d�ZAVV۾�WD��M���x�'m$�(O9lC�	I$����FfO�K3R��9�ۢ��e*��6WgV)��ح���	��t���G9�V�����8=��U�OK�]]n���>�3͞�n A�s�p��3s�x��v�V減cé����Qz�;��8P{]�o�f���Y�{qh���[�k]Yg��Y]c���w=�s���/<��ݮ]����C��ݍ�k���'b6�pfP�������J���T�����z��;�vb��ݥ]X��p�eI%����P�Y�b�&Je�v�v��
1��D���FTA��W�/,,�fH���mxq�W��E�$�bƊ!L (�3�Ud�*�x���>~��d �!�Lb���
��Us�d�7Eh{�}sE,�F��Lq��G,���_��W����m���Q ����h~�J{� `~�0��#�-�f�x�tB&$H�l ���|���/�~����~�ʬ}��?р~����~|�ѩ"��\���lk� � ���$�$�$l�$pƫ��?M�>q�KЃ�7x�%��0O�߫���g�o����%�8n��*/&�I���o��?{�����f���{�~[U_���?�(��!����xmm��TTM�O̘�_��}m�����8u������5;z�ٶ����w`Z0�_�Q�b�} yx�rH�	�7m�]V���q��'DdQ@���/NO����H/��gR��l��� ~���x?X���?�J&�H\2<����c��0�[��.��1�j����}�+uIw�b���/�E�8�r�ьS�ۯ�⬺��f�X@F$��]�/-��A$���A7!�%`��=�p���7^{��o~u�hIș�����M���-�V}X|I#�,���/_R]�&���}z�f+�Sj4�)H؀��<58#�2�y/�oOh�}��櫆�1)F�U�h ���$^f%Q�]l.1)P��?@�]�)^ ;Δ�M~P�?�A؉��N��Z?*7��2�$�I%q�K=_g�����4k ��¢��ۧ7N�Q�2v:f��������Տ��C0����p{�x�7�J2�5�!��U���"U��%�6���qѪ,s�u�4|=�7��/���2�8�d�$2K�1i����J��o^AP�������H���X�HM'���(��A�� �c#=!������n�����8�ˑ�xSy����O�b���5�A�����b�QR9{I5�U�*QU�Ȭ�
EɔI��*rr�ř-���p��_�?�J�޸7oL�o�x��k ��߽�1Ş�c(��w���k�� �@��%����.6�hm�F��L��٤>�f���7���]�u���MYl������ͽO�T�ۼ���x�����˺�ͬ���b}�3���H*[�+�:>�Y��#t#�8��F��͛���(��o<�~���dmW�����֙��z
��e���;�8���A2�dD��ߵ(+,,�F$Eb�^+b�"�bE  1<\�(
H�a�:���X��]F7߹�4�!����U]� ���8,Qp��Xt}"w*�Q�IٖM�?@���|WyϠ2�"5��Q]�G�|2�n���gd�[9{�S�5Ʊ��MC��~�|Q^����|Nh�:�K>�|���v����X
"����%¨��gf܈�!L"�^��+������Ty��0(���s��ʛ�v����Jx�1AE}	��A�q�eG�;�D�,�2��24$)K�张J!J���~�U��i?�X'"�vL:��eh����{���xQ���J7H8�v�AS�)�y�m|���{3>�K�׃~��
��\�r�N�d�_;w�_@7!��b�	(���>�O�0�SBW	�Wμ�eּ;���7�g�9��p"t`�C�m�����0�m��]4F��u�����~~[i��%�
VUG�"�@$�ON����c�%Q�j�����Mjʮ	S�|V=Ʃ`��VI6N������H��܆+��a߳����㍚Qk�]ڕ
�2~������a}_�����>��$���UIex�����uA��
^VWhW׎!���T5!��>Y����6]�������	��O�$��O�K���#4v��u@1\����L��s��*-Ov��zY
B܅��Zi|=����| �|`x��8��*�DC}={���U��FR��,�h�Dy���9)�<8���,����A�4�� �V_���)����ӽ��}�[]'P�#�����u�����/=�\kp�^�Iʋ�t�T�9�;I���6z���v��^ݵ�����:�v�	��7e�����l�#2G=on#��v6S'c�yn�c\�����^]v��v�N{Z�⛲��F���f�$��+֤���
�-鍑���Α�æ;:�v�x����*z�e�����{tǎ� ���
1�� ��}+?Ht�*���y�A�r���]Z:X4��I[���P�q\m�^z�ꭈ^`۵ɨ.6�[���fS^��0Z�K)�$��m�Q�C>�ȋ���>!>�p�Q�~���;q�S��Q��a��I��m�Ô��?x��(����=Um���d+��/Ԇ�D�������m�b́��������`fHI
f���Ǎ`��A"�DZ"��c���'F����C4	�����\~q|���%����&"���-S4����{��SHv����<=��!����o�/�+^�\��A$i0\
�)���Ć��=�pa��c��^f�^V�u�-��F0�A*��$��RJ��&�������UUF
��X|��,`�
��k�Gu�ʉLnM·���y݇�j{q�bkg���Ѯaa(��8��� m�"I3�B��b��Gk1�Ty��Ħ���Ukw�;��/1�� $E�Ϥ%�p&���lƤ��%TLB{J!wߎ��᢮�~F��rAfZ�	�\qfEC�b*��5b3IME0�*��N4�1��"�9%�����'���u����K�?�򣹱e�t'�p���:��n���������IF9�5 > �:��~NXH`���2.}�8�1Vj�����.�I�'����+ߚO[?�����6;�}�{���~	`oO��e9���F�|�kW�3]ۛ��>@R*��;&<�NO�{}��<��+\)����ٔy�����9TE}޾l_��oYmE�@TKG8�]�u��S�HEPRZ|g���7g�߮�Y$>���e�&���$N�����Ҷ��q�G=�\S���wg��Jʜ��w��߀]�ق2ӂʉR|����B��tsCY4׺��5�= ���S������
��$)9�:'�!������;�Yך> oJ���Tъ�9�����i��Q ��Y �RNF�n��b�� ƤUD8T�C�8�
��c�d,�
*����2�75�VC�����cmC/q+!<r���_l�w�=��p�ZOeb'_w>J�6�塹���^8�$X�ǲD�S���HP��wvM�P829G�Y�MC5nQ��H�A�\p�.!�u�Jޤ�h��Y��1CX3��H�^<9V���0ݩڤ�F��|M{�c@�ш�'O�8XU���i|v��V�/��wCWw0�Y#Я�f��w�q·�I68��ʫ��0U��tQ�K�zl#��-��J��2i��tks{�c��)�����ܱxD���U�p^*�j9M(>��,�!�t��U�ϝO����OP����_ܾ���ZF3�n��l��Ŋ*��9x,_.�}�nыT7�r�eA�a+Jq�t��^FR�VW�/hCk�de�vx�K��]:4G��y7i?}��e�R�0���t(G��+?G�(�dj�R���&��u��B����F212��C��o%ԵWz4�RѨ�KL�칹�[2Ĥ��ha/��l�im��Pݪi�0��� Hay�
�S�@Ϩ�i�t�Ȟx٧I5˰��[V�:�r��;̭�I�4K۫����`a���4��^�Tƫn�G�ח:��|{1�b_U�w4�<�wj&~߃y��3+��� ��!�y��'�W��2��������EW*�k��O$	��n��=UO-DN�(�Q�z��G4ϣU�5y�j�Щ�8�j�y(cN��d�m�~�&������n�\��>�+6����iutݹ��j�W��Cee��j�3v��,tf������E��!�ai˙;�c4��b��[���ɑή�1��cl����4��~�b�|�u����H�
��Y'pu*Żk�V��VzާW�M�h阻s��k�Q2t��C��B�,����u��LX�8Χ�mr}[��4^m��������PYm�ʕ�[t�ͳG[t1�-�l[�SJw�����Qe
�F�c���V94���%�z�fvں��̹:!T�r�jn�U���+d�^ʅ\���[,.�Ii!s$ʌ���k_��0!����0~"��ߛ��j@�r����:��Nٌ|G� =�=�Z?/V�����pX+:������c����B��7�0\n�7��`�/,P�d&�Q�c���=uӜ�$��٢�VM5��^:��ޅ4h�*	$�ϯW|y�~�E���1H����wg#�!��qX�0ej��79�Ng��fۆ�q��st�9 {����~�u�*#)z>��|�<�n)���m~~�y��(>��������(8�dH������P�\�^������j�G����~�n��k�"+�ܹ8x{�}��1)
�$+THb�?O�z2��kf�>����$N��wzN�}"�ဌԇ��d6��� �Z�1��I�c��c��Z{�U_���n/ɣ���N�O�:��������܋>ۣ=�贬��ڭө��;6G�l���Lq"	�������������IX
��s~�\�]dI�-Ƥ�(D׋qMh���N&�ϯ��c���o��������?�(��O]����W����nͰf�^Ů��蛑CN���/���Me�"�7��
2�Q�1����S��s��9o�񍒢1���_�����m�F!��G�z���o���8�L�����~)S�Lm4�ڪ���#��X���%$!��sM�������BR�A��D�K��>�>���KG�Ls���_(�_�^��ి<=���jl�F�Q5da��~��?;&��_i"�������w�_��g�������1���o��_/��<��|��J��s�18�J��Q���#$�F,�h�d".R�G�ןUQ�5�q�e�w�}U���?�y%q\�A�#l%�Wl����O"���}��f\�QO�ۮrdu
�⪣哇��*���'���U<���;��m����|��+���u��T�nm�/s��m #$�7QƜgq�X�+��<MIė=X��o<]7H�ټk.�l���g�t;�pEmy�=���Ӵ��&4��]������3��z9	v�ZB��g����[e��k֗�6+�m۹�Nz����\¼�m1��m�F��n�:��n=]=v��MΊ�z��N�ɞJ9��1"��8��>���+�^I.���d��*N}��[��P��H$�5L��rmնȄ]�z Ֆ$v랩��{[�c�svۚ�sc<�Hp�A�x5x?3��c����ϡN/���|�O}�q�>��w� ����;���� |/eWO��YǱ�՛�+�ƹ�]{�X#������n�Q�������^�>e��X��:���p���o�U,(�H�62?x��ƅ����ɄtT���l�����~Lӈ`��#~\>���z���lW����Ǖsu��=���>����ፖJh໼Ul=����"U�D��������w׫�����9J�َi�V��U6� ����P���|��R!�	�i�J������v�۳{8�ZzWXn�,��槾߭{�~?��LȜ�x�	�^w���>�H �O�0M���!#���� ��\u�x�}�e��0��0I^���M�ߟ������u��4�$�g)�n��-#\�[��k8�<	�n���bW��^�B�e�{�r�l�r�:�QΫo>;�w���|�,QH�:��6�;�Y���;S�kXcqFhAN�������lq&u�ǫ����y�I}uF�>� 1�H�}T���=���ʀ�$�KMR����z�02�%k}��c'�c��*0U���E�J�q�`�h����>�{F#Q��?|��b�N@����+�R�}���GG]qx!�����w���i7�sl�ձ���la0=s�ͨڶg=n�����t"^�����IB���u��,B�.�T1gX������4;�>���]_�k���V!;F� 4_�0�(c(�Ԫ(����|H�BUi,���@�Ƞ1�$�ID)�e׺WC�@&�ڷE7��C.FS�"�&'u�sG�x>�U�'9�:�~��Ļo��nŋ���R˭>�S�o6���k^^	Է�n�'�C����s�0���(D�������?�&�H�uΟ]w�ѳÏ�[>�߸�4:0��T�UG�S�|v�9w�O )�3 )�*�*lw��������ش&����)�%���-?Sx;�������*�*�}G������ps�6�A�燮�V�pدp��@qݝ��r?Ϟ߷���ȦR���A����R���2�����jO�L׿_�S�hG�8����T���WY�o�d�j�����q�s�"�DfzgK������w��^)��{�u��m�ſ�B|����)8�f	&_�#zSB�pjBQ�Eޗ]��	���{r>�GTb޲?�a	�Lw*�����t8�B[�9���������=j?����Q��Q�5��r��E&�r�P�M9ː3�ې-�W�L�58��*����*�!�}\H&LQdO�Nb����ͩ-���UQT���]3Ooy׹|ti�3����ӱ��;Ecl����a���'�ãnEa2����mf�a���:\�ө���]c;:]������?����������uрܱ��73ƪۓ=b�Q�)�N���u�3�l/c[�������Z��*H��!�g�ְ s/C�~�4����U���3P���fC1e�v��9���a��au�d=߫��nM��v��Ǜ3tgbxQ�ڏ��~.�$Lp�dq��0��(�>�O
59�i=����_��Y��W3b��z��!!H�R�H���מ��n�y�n���Y�ՙ�0L F1ȉ�ϝn�"bI'��g��$%r^?l��"p	��I��CW���u���V��0N������}FO�I[�ZGU[�k�����#�_�����U��om3]u�)�۶�\��um��zl8��:��#0�]۱��t�[��9�b� ���GL��;g�c��\�I��ƶ�]���.*$ݚ�{cհ�4Wn\�5mݮ�ns�#�Z��zJ9�u�c�\nuq�C��\�`3�u��=���p���\Xݞ��"��Bk�EoF��h�q�p�%�˗�џ*��pj}n|cfP&"O� \%�_��?e�90���9+I��l�p�������Y!*������cr	��J'����b-�;Y���WXA�׺ݱ�G
��nV�o�����TZd0{~I����Gi��Y��l����j�(HXa�B���� Ql�>׊�\��`�z�����fr` ����Dh�h�q8�f8�I��Ť�Zw���B@�u��V�{]���N1$Qa�,h�A{���.�)�0���-��PEЄ) �R4{�/D6f���)$D�;E{<6s�dq֨�U�xM8�*6,��W�|�+�tO��D��w�]g"�F
�$D���/EG����:��U���gjK�1D��6X䮧ͺ����@J�7�&�+�c[�=5R�͗f��.$.��������ߊBc�=�a����CIA0j�N���Q�Q��R���#x�B�W�ߒDr`��pʹ��9ĕ�L9dX�8&?�G�=��$�'N,�	?V|*���B�Q�����[�;(��b��K2$BZ����o�p�]��)�&T6K�$���o�{��|h���Ǒ��gY�B�~����g�m��b�):�K�h�_�_ǠQD\�&;ƯPy��1�E@`,<d �=:�Q�gA�����X�M��>X>~\˅"ɒ�:q�%��f�C�vWu��a�/�5pF�E��Il'���}���3��P�P��.�������pvMv������9z����|}�M�%��,� 0v����k|߻��w�Z:v�V��%�5���� ���W�Y�~���wx{u�n8�������wZ�â5<I�C�#3�"a	ޅ찕�3[|�A7����23w|GH�W~��T��tc���ʢ%JR�0"���CW�"��N"�Ä�K
��Ц������7�H,���8}�m�|,�큭�C1W���g]pT��,ݵ�п~�R��R�2�	��G%7Bz���##4�YKSA��tR�����D�j�M	'��!p%i�*�I��DQ(*׸7�F��a�0�i9���i!�L?��|�Ƽep��q�1� ��h��5Q1A�؅���L�b��ݻӱ��[�g�2aD�	�Hcj���;=W�^޳�&� S]J���t��k�>�\���Cn�|�4���E���B��u�Dd* 2S��C���=�D K�c>���6*Y.+ADDl����U8�6��[0�}��Α@��_)��h@��k�(C����S�C�2Zm���r�o!�:��ŀ�X(�2�̩VB1EG�U:�s����9���oej��2M!+�(�І���g��q�0A�X��6k�cW�3T �J�t����6�JCuN����=���/��@1_���c�sۑ}W�&IM���[u�S=Yj��T9�s��k�cf��e0��y(r�o�����k��h��׊����9]=U�����Ƀ�ℛQc%֪���QG=:s<��{�z�D�q��
b{O�sHc�&������He���au��{��GQ��ґ��l��(?��0��	d�x-��}4���.�I�>{B$h6-�=dEEB��]A\a �@$���fEIQ����t��0`�Ɍ���|���5�}��ֵ���~g��i��>�K�>3�,���9R]%�z�V�DP�,�?[����#B{H�9o�>֍�Ȧ��zsI����%�ƿB����*/�z�-}79��9	�G�#��P���ӍL�t�VhQT�7H��$ƙ��2ma��w��M���>�&_���,}o^�������$�o��Z}y�/��������Q��	J})vؚ.ւ0�}^ڕ[A�v�gț[CI�[����_qc+VЗvҮ��5UeU����!�uت&�!_GV�C;�N;z��UB�$�_���#�|/�q��W��Ɠ���}rJ�q+Ds���9���e^��?��O���b��~?��������":�m1񏙥g��C�����1
���n��S�iԘ��:-���4���/Q}���w6�ز���������.|ɟVU�(��r�5�x!)ZA��C�����:n��p���ɹ�������,|��\i������8W�*�hӅ��uf�W�n����X��Y8*��U�O�\��?��g�1�Ry)�-!�����-�ޠc{��e��mz���Y���?�)# ����#s�]S&,��
c*��ž.�j��߭�Ɂ��^4K/�`�#3�uS��Y�]Bº%{W,�vbe�Q;k�{�7u�;gm�[m��i���9�K�_�n�Hs���3�`+=,4R��[�v���N��Q#��6OELp�/�i�S��!˯j߯V��~��`����[�ۧ?f���1�I��=������NUIm�@R]�Y�ow%�wE��I0�,��/8@�ŕ����A��Rr�4�;[�B�G|��3��kEz���{T���=m:�]��n�*uz�:G��T�7�d�^��O�ۉ�?db�A�K߸�!�*��+ �̀��g��uzT��j����Y����-��@�>W��3JM}��L֞��\�9�B#A��u��B�9�}�~�>a��u�L=�ͅ�vz����<C��W;�ז�/@�ǍI��m����؆�ZȦ#�vۍ�
�{��v܈�m4,�g�'�t�r�1�n嚝=�f�V��2��r�1�g�q����g��ۤ�q���7�ȡ���aSk��n���:q���!���@��=��%�n8�tuqj�W&;<���]3�<a	�qd�^W�c�41�y���.�$�w=��øgqA��FH��w����v�.(��prC�v��9eS���G�plu�փ��-�w���+�Wr=��'k:l�+s�OӰ�r���{]v4�w���un�0'�;]N���_��|���n���xKgq��ͭ��]s�s���I����{�#��#��Ht0��ݍY���;�q�#��Tr������1s�\\�e�\�qi�Պ���	� w�b�a�e�E���q�uʻ�mn���#�����۩GD�iѥ��]�ů��t%�9�x�;��9I��r����nlr-�3��b�v�e��nz��.�kwGQV��X|j�o4����u�[g����:�=�v�Bq�y2�=3���x��Gn^ݍ��NC�'�ݧ�V6=rY��u�9�On\:�Y���S�޹Zn�ӱj�j<�k��Rw�y�:=n�J'pH��
2��=]��WlI8�1��Ʌ�����rc�<�vM{v�a��6�#yR.26���g��llMv:�����ԧo6���-���r�e5s�#=o+�lM���n�uTl���.�^_l��d��nNGM��Y�q�u<e�<su�ېz�l���\d�Wu�y^�x:�n�X��=�q�����ŵmE1�Jض�\�[v�bק&�h�r����Z6�n�Ւ�6{\�,>'t��ghh�v�:��-=n7]�6�6���܊����[u��t�W�	�۶贋u<z�	-���F2��ךC\$��ǎ7��F�<�[�]k\�І��[v(:�pE������g�3���nlޛ2+J�^�i͊u�[�6��L�@��zC�c���w׬�/��JxvywF�������\u�����u�6�V[/�ޕd���5"N9��od�T���S�}YEmCd��ͮ|�5�V������ ��s��sh���]�gn��!�kF��8�L�H�꺳re棒��[�\%m��e��EɚpM��ga.d�&��ʽ����]u��X�o �����S�g��h��]�Ζa'�Ü[�:�r�2-=��T��{5T�
Aw�Z�V[r)���oi;JUS<��;�٭F]()]K0��3��b9^S���i�P�D<Ƨ�q���ŋ�2Wݓ�6�ڝ��Ρf�V5�S�	�EWS�㛧{��r��y�ؠ�:.�l�qX�b�Zܷe6�Y��w5*j�mR;�'Ml��^F�g-���Λ�n�ڝ�����j�Om�H볲�#�v�r�FtGj���e{L��7)�{�]���[����z7=��2�>���R%[�
lQ�X�������C{Vz��)K�P�\F�L�I�K�G�������}�[h뎺N��Ք���(���G��Wa��i�p��
g����0���s��1���H,�H����Uo�5������%�Ｒ�Q([D�ʤ�
�l[�)��k�xP�\�{�G6�壧ȯ��ߘ�O��d)�HRZ�H~��@]���� �bVL-�Q1k�Vj"AKi�b�oFy��q��b���׎-�oY���QsqQIW�>�����(|1	��`�
�+�m�PE1#�.\N!j�߯8��"AEUR���
xQ���j�c7_͋8��4�}c:�9t�hَ�W=�t�n��p9���9��'e�K���HNv�����_}��;�W��1�R1�SA��su�T�s�����P�;�ƾN�&�LVs���w���X�X��
�S:�d%�F��B�r*b$a�&�(�h�D�TR�Jb�$�哷�?4A~ �H��S#������w��+���ǒ��=�+��`���p]f���pxxg��s�����j��/��0��8R/�H!����"�7���:�;�3�#DII�A@b"������\���lL��Sb�#�#�⨗���<�|����̄K;B֜��ݍ/��(����dC�3僘�L��lmò�r$�"���!w*p#낺�_}��}�7\"1~:Z����ㄒ��d���+�ۊ��}�:����b�mY6ٲ@�s7j�Uˏ
��i8R%�a�.��ץ5iX�#,a�W��+��.z	��r��~=CX�7�J*D�M⋩�lC�(��kO�!@�`�}� ���7���"�+>r��U�2`�b�"�VTL>��ܽSy�C\��u↢P��ѻ�qqU�Uq�V�n��A_��{	��}g��ׂ�@�?T���Q7�)v��۳7�Y��c�Q"��@���Ih��M޻T�S��a7q/�m����!^�p�Ԑ"��;�/��������	vm7š#6�qBgٚ<]$E��Y�����:/��q�˓]|�.5�ލ�v귚�6=��X�gLQ�q�E�0(�8AųӼ+�����7��@ɽws��y��x"8�
)�B`��~hM� ���W���9�r��(�7�~���0T�ƾC�huU|�p�I�����l�э�x#������p�n[
�!FA�8c"H!�������3ԗ? �IckA��Ϯ{����U�m)��z�X�AӸ��0������"d�����߅)N���A�gV9M����9�����-U �NX�HIe��K�5#b�,��.L���|d�s����ċ��~�{���x�Ǻ7Vf�w:�N�\!�;O�����M~< �O��C��R8�Sɗn`#���O\^�������8q��Ndy	��Dq�N�n����vNŷ8��7m��筌���'YJ�s�tVuH�¬��k�n������
B~���=�j��%��cXg$,��]3PzL_!����4 �1�Y��A}�C�c)��?����p�f=o�CV6��ܺ�����bFQ���GCx}^�����{�WK�1��	E��E�R^~��ˁ�^hP�w���8_�A��j�}p��/倓�"v���yx�{��E��O�@�f&�R5JQ��P�=8�
�ϩ�_Ԝ�7��^��֗)��T�(,H`��
�o��Bv��I��N$�Y�/M�.$Ϩ��<��l�3�ے:���4ML��7��K�ƣXn�:!�V���(r�&�z�R7B�i�f�z%��냊Y�k���؋jn�v�2�!�Ij���=Q�-ƀ絹�n��k�-��k�������U�໵ݸ�UӴc���-�A�v�-�M��z:y������>ۮ�/k���-;q�F��1p�ѐ�7<�b;v������;�\0v�[�b��`��vx���\u��uQ'��Q�߾]_�����q%-4�,�+/�	�!y�M��3D��n���պ��Ƹ
2�cH�����9�KPy��!ͫ4R�y6�]�Q�H! ��	��hW��<� ���4��ha��}V~�0{l#_9ك�)��,�����B�/ 4�9��(bF��y�~h>g��d�C�Ua(ڑ��
��ӌ�^��Z���XőQ���6��Mη���u�1%2�F�e���X#�&;^�1���J�m[��c�A��Gȍ��SAU�M��>��Q˛Cw���&�b\U�đ9��׸d<��ߖ���̚�"��N�������("��?=�Ux�gp�қ��FQ�ڏ>�~����I�7V�臷SM�cG5��˹'T�����c�����IK5�Ե�3�"�.@AF�AŬ���i�Z�D
�y��T"�����}�ޅ3��SSU�@�3�A���>��{�5�~�?����),Z8�#!�Y-i�/��ˣ9�J���.��i:ϥ
�F|�d�*Ӓ�
�t�`8�)"���{�[��`���U��R)��LcE=�SF�1��n�eG}�͆�6�r5-��ACv�5��jOf
;(��ŧS��|/�)��	����ȒR2T�U_��b��x�@�?��q��-�X�l�+�P �RX �,l��r�;T
�CxH�l4B	'��
QB�"Gg�6[��<s�e�#m�c-���2���2ڱ���H��G"�������w���!�۬��_e}�R���{)��M��B
(�j%r떒4��4�E�u�}A�S���`�PQdUQ I �����}���p��N�۹0 �sgy�]���w�g��F*⟕��R����� ��(h�*�8U$��%X��E��I|C �
O�ح�]�Y��
˻�����]V�_]��fic��xg�~צ��5�,���I����6#q0�ͰC���:��X�`��Ø�
z�j]2�²A6��X X�_6�h����\H�kټ>���c~?}F�uy��!�(�-�[��2-�,��_{J� B2��24�y�d�umH;YS[���Ulj۴=pge�|�{>�}��m�v�9OH܅��|��X���8ņz�{�=���E�P�R��m�9��&�A�
�!�Y$�͓b��������hG�!�UQ�"1�M��0L�tۉ	5"�ۑ��#N9$��.:
!>����>�<���ݢ*�-x�oL>�:�b4�-�*�HC��]�p@�e���4=�=w܊���,:����G�Sa	���E�(��9��p$�f�U��h�9MS���`nO�IH䫖´?��B�YU�
A�hH��{���	�K�����
{�#C�u��`�=���ָ��i�̼���Z��ӑ��M �e^py0X�E$�� b�3s�/���DS3Gts��:���B�p�0�r%,����v
hHʜrw��k����x���]B�X�3I6����TSH�*Id�� �#i�Z�v��Q�H��<c?4�|��7Aa�P뙹���7w�����2H��H�����H�ۯ��u)��(��F������l.Ĥ�+��ฉ&4
F@Z,����ג�Up��f������7A��j�sh��ׂ��x�#DO��Tc���)e�3}����j4"�6DB�DeJ�)��_-�~I�)/���9�;����qOR�v��R��(�S�������Î6^X�8���ۅ�X�'��.ݺl��C��히����rn.w\�v��Ҵ�ް;o"*\�BN7���l�DwlmĊR�ڴk��1�=<��+�ϰ���/nڣ���n�v�������b.�^�}E���<i8g�cd�+�h����H	Q�)���ɰp�4\�{k7l#��Ϧ�JҌ�\��d�Rz���h�[��eFD?]F�m�v_K<�0lGI븽�藓݈Bs���X�Q�;Vݖ�<���5��d���:޿7��t���t2����ص؀Պh|��|Y��@�=q�X�|�9!�E�BȑpKK�n{e�#O%{��䅁�$կ�_9߄���}��>'�|NY4�P��֝�L�u|�A�p���-`�o�D'�p��>��D@{��wo�7n��=�i��3q�$�uᚰa��/c�kۋP�o2sy6q���Ƥ����1WBAT;���R�/3��o�(��C��s(�,_���J�,�Pn7oP�W:�W-#Z�٠��=����gj���v�_Q-B��ƓD8�\�8����F�`��,<�����*^�F|�q��q�w%�]P8�z��W�ԅq*D�!+%�K�,�$i�P�&C�ff,�	??�r�_5K7���]x�'�ht+���륓3��~|}��o�EEXb
(ȴ Jm��/>�rkʄ�lV#X��-����<uB�f0�a��a�*���G\�	X�~S>�x��� f��)0c6ڌ���nR���Kg����J�-����ߴw��W���T�ARI F���Z{�JX �(��S�w�,��0���+�}P&�W����,eq������mġl?!#���3`v^���^���n8}���W��"���������3��8\j	a|Z�����f�N�ѻ�G��d����{�c���l�Ғ�_do��"�4�A>FTs���c�gB��(D�A�"��@y@�O_�����Ew���y��\D��T�������ܻZ��5��~'�
!����k1[�QX� QFIV���*�Rn�w�R�ظ��E�&ZWi*w*�fY���ym����F��>l"�䔳S��qr�TH���ZE,EiFĭ�PFi�An2�'�)M����CƔ���5�L8��nSٓB��*kl-�ӻ��/mAf�^k���,�m�(�0$��#��FŊ!����ufe�:���k3%�1}'U�s��ѯ;璘�{e�R�P�R6���W��KE����Eu����E�J���uҞ�3��O4~l:KtU��ܱ��쬇�D� ��?L�9��I��L5
@|D*�&`�C깸�����]�>�	�T��Lߛ��`���Eu�$.��D���~�ϲ�ҿ�l>5���G��vĬ�+(�֯b�B�����P����X�gi�f�t�DX@� �ž]��;�%����F�Y[�P�t�:޼-�!�PB·5yS�� ���W^��_k�ģ�X�+�j�o��AX��F��2�d|I��M��e�M�m�+I))!��k�G�Eψz�;����M�9$�a�(-y���-2L�@ZC�i���#�l�y�ƅRY[�Y�>V)��Wgۿ�U���c�F[�̻�"t����haM�����#TE�J��CD��PZ��_��b
J�!�.	������ߛ𥳐P�IQd��_ƾ?V����h���le��gI�mD�L5#���jv����Q�V��/ګ�6�v,��XJ�/���]���+5��F����ꋰ���5P���/���]K�ո��n�^$�F�*�\i�]�k�Nk�!ҩZk|b��*�:�n�؜ĩ*�e��֞����W�̝.�5�[��X��@�^��ʅ_J�"���ݧ�Y�����X�5+���C�]j��:��C���,�$g-�F��gS�R�a��9Y�k�ܰ�`��.��n=�]yR��w]��C7b����8�ۖ�kxڼ��v�2'Q�ή�����zY�4˙�M6lg�ϒ�s��]#�9q�����}-K�#dw҈����/��Cp�<�u�U����<�b�S��!��|��fQ};�H}��_��ߏ%��/�IoĖ[O�F�:y�7rZh�J\Q�"����$���&ʁ�g2�0oT ��b8���}�I {��V��Y���t|�;O��aO����ɧn9!0��FQ�'h��� ���-�lY1�66��M?���^�����"C���p��l-��S�nCPHCQ���.ϖ�b���ݎ@�B�����3�(�pfiPq0�d�Ɣa2��+�m�`��-h�6o��]�|�UQT�UL*g$�Iefkh���rT���r"ʚh*�E[�8�Т�\]ܾWCdK7�X�����Nݻy����������\0�@AV+��@>��s5�,�m �H���Z9�#��	;�4h��E�|����m)��F�l������Iy-��:x'���	&#�$Qbf�R��@�D�䈘=Pv��?x=���7񋰜;G�7�����9�� H�E�{��7H���7$���Y���"%hlA$���o���f��O^�Dk�X ����#0���E���>����4l�D{N�pa�/eZ�"�i%�D��-� �7��+us\�ʸcVd�4E�E`)N�VLU�kuǏ�S)��,�	fBȽ���>�]����3�^�v�
���}�t%!'n�^��vl���y�]���8��K�h�%d�\C�$n�՛(
���o��`��7	G=�9ֳV���щ�x�yۋ��g���Kd�n{c�y2���'�k=�;	����c٭�Y�6�9�����[�u���� �M�xm��E�K������8R�R��sD��w:���W���vդݹK����a�g��r]#ɲ���ۭڄ�k�_<���S�#�F�v���1�L��ݗr �0�C��I�$�#�+�(G���)��khIF����T.�5^\����1����qv$�'���sj�Mqnz�ܳpZ�I!�;hl��=�h�I.J4?_��Z��ټ���F��.��}1b{���Q�m��D�I�ܷ�J���eQ4jN>\���u��ck������Â��௾�K(fx�x3��
I3#q)$�-�[�C8|#ē�A>�:{�Ck���(�=��|.����A1M�3�E��]E]���k��{*�r"(�{)��E��N�e%$I�#q�X,�����3�R� ���m������w�!f�����cm��;=�m�cU���c67qv<=r��k�q���]G��j�zc*��q�Kw�,��,h�:�������0��R$�$��g� I���}�����%�%pq��D)�@>����'���o)CtiĢ��⨧yڣ�igZ3�ky�P�~Ե���y��w�,o}mX� nB�e���ﵭ��jҢ/0N���dئ�p��Q/�t5�Ȣ0B�AF�$�}����
ٷF�lE��*�H�UUw���]��l��qT���WGa��bH�0K]��|%���]�����텑K���Ep�x�c������G2r��.�X�=v�u�۔��G�$�#AHIV5W�bA�@�e0Ғ"�; ��N����gp��ȃ��[W��^/�R1e(����A"��3�#����T�Fڐ�Pj7�o���Jh�)�Z�G�g�o;�j�Bpf�x�_E�2I}Z8~�����0�B}��=��:�u����J "��L0�8����(.H�3U��KY#�dT*(V*�H�����U��O�{�CD&I��~5��>ƥc�v�Ű�g"���:p���
�;��'�4�E�]lc�0�=�8��$PQa5�v����W�7�7G}�Ҟ�q(�0��P�.��_������^���
����ޅ��k��H�����͊�v�G����`Қ�OXeZ�'Wj���2�e��"o�拇���u�i����)��� {s��x�I'ؒ(�'����{��w�{�� �(D� ɴ�Qұ��2�e��e��a��a��7����o�H�C/�?F֍������L���hD+���;�!�^��w���l^���__�C�c^h�F�"6c)��Vn]Wő���|��GEA�i[8�?ߣW���Ȝ����iX(�8rn�q���Ɲ�j+��K��l~�YV�!���<��'���|f}�8 P�"(>�Gw�
�+a�I[�^{��8���C��v�ȕ�Xbf9l��n��,'Eګ�3��Д�/ u�5�j�������J3rA�%��6=a�0fhV�[��2�ғH�m�,'�ε��sq�bƮ�^���8��te4�)����
�Q���dT�V�C/��sJ?{3~5:�pw��ڎ	9,�M������9�װuQ���������;�b)�cPڞ7g<��с�C�_����^���P�j''2���i�ӽr4$�B�r�mX[�-Š>�E_���d]�V�tT��F�ǩl#>L�\V�EI�Rx�uUdY�������Òj��0v�uIv�;9붼2���޼tu�J��+��g��$#{]�X�9��6'���t>zWs*�OH�r9������v���s���㹩ã�nxxct�.۱���"��b���q�wmᨮ. {v���t��-�v��� ������ts�Y�5��]�s�{^�w= x�u�l�
��%�,c�~C�L"�+�L�顿:����a�.)M��QF���k�7#JF0�����zq���{1�%"n)��>�b3���߯��`�TJ6bD�S����F
g�c{�&j��D�V:��r�ڊ�"*�*9��G�{;�֨�������F�PJ1�q�����o>��`ɜV����{9tnE��6�(l��YL"nD܈�����2`w�=�C-1sh�|��� |> �<Z�&(7�9@�y�	�}�~7{�W
^܋��O]F�߹�j%$J Ċ8�(�߱��.��>��։8f;��3E�F��iB�#�u�(���.�]����.�wc�;��v�GG���t��(��0b�u���՜�;u�0�"��AARN���;�bZ���yp���z4�_-vtH�#f(#%$�"��/��_"?%#D�����9���ęR�EEEPU�r�Y$pJlY�]&+	�(��EG�n@��DH">6��!v~��j��!Q_C(�l꒥$���f���O�*yXH����Z����ﾥB�0Qo���)!���]�����;_�������<|||����������g%9Q�"t�#�t�p��>�ྸ3���s��:-`C!#4�M&C)��b+,xߒ/׳>�h�oh�8���9����Z�*t�vd�Bu��rS��Yu��Fg����~a��r#�|�Ԃ7H\pF���w'K&�DW�;U���=��	�b��Q{�ϱ¯E=�>�_F��325,k��O1!���%�Y�Q[��`���S&��'!n(�?4n�^;ƳK#0~����FT-R��U9.6J�S*��!L�*��}u��Y �3�����}�F�=Ĭ|k;��ztf���\�r�қ>����X�ʱ�]�Cl�E3� #����C�v�=ܐ��ֵ�yՏ-��Sȡ�����5m�"2D���>�H�����!+D�ƕ�|7V�^�ޅ>� �H(8fJ�(Hb����[�����qmμ=�:㷱[e�W�+\v�L�Nd;GX���k���	Dh�]�&I
iC�8��ݪ��Y#�� ,���r����Ш*��3?jޑ&�iC"N"��{w��Sm�n�uZ/{���Y����:e��8.q'�;��p9�&cs�4`��s��h7����"ŀ*$���b�{���U5����REJ����kꦧ���pr����<=|��43ฏ�~���.�d�T���:�u��f�e<�G~�ĸp-8���9"��w�W=����ˣ�=ݛy���H��TRu!I۷Cۮ=����4�D���D�/:,2���6��܎��7���^5M���o��6.���^׍wv��zLGSX�PX*Ȫ#6c������|;��G��-���ŧvy	#�����2������Ǝ�Gy�ŀػZ�Vc�d�F���f"��w>)
b�x��^�x �D��}�{�����f���o	Q� &8ԅ�q�U��|UB�}>�7>$��������M�C��Dw��(MH��!�sC/,��j�{�$�����_�s����H�9�굄��n��*�=��ADUЌ�5kR�@U�@V��j�	�] 	W� � *c1�.��1RZ���
�=�Pd R�#Dj�*RkR BJ1���Q@�Puە�j���<�0DU��s���4�-y��A�U�D��G�����B&�9��w���o����{F���=O�3M���Mi�U�E^�;;�8���Au��TEX���Ó���!7��l�� ��6:1����xw�Z�c��E^�=N/���¾I�S�����8:�0���Ģ���Z~���~.�0�\P�yN or�̘�_��/����
���� DC2E�L�Rdԉba3�&m̘iɃF)(#	������$Y� єe	!fX�F�I�	���	HA&a	��M�ɦE���l�B(�L�%!&��2$)J ����d�&����!�I�,aF(ĉ�dY�ѓ3I"b�F(�Bb	I	2��B1D%2��b(�F�$,��230�H�0̛M%FK	&M��	3!HEF
�0E��L�"�D�2RRHY(2&IS1�bh Ĕc�$�	�!)(��4dH$d���Id�+(��(d$�2Q&C
A&	)��$��!��0�`�&�"L�
(���&I	��	�1Hf		%�I	"d2HȒR�Q`�3"AHAI(d�&&Ȓ�Q�L%D�#f$�(ŃF4Ča�JB	$(�d�C($0̐�1��6E �d2L��d$ȘI0�)��$ ���I	�1%I0�%�"���H�RD�3	C#2AFC2L)I	1&�#4���aLĉ"CeI��f���RI���	�"f�4$d�%�)E���)	��!!M��2i��2bMD�4�D̔dƙ%1$Lh&))����I1�FI`� �&fh��(��d�)&)!����2MJ2#IBh�#d��d�LJD�$�Jef)1d�3J*E,Y4Y4i5�f��i(�b�J2Q�J)(�F�%%�M�M�M,Rh��Y(�Qd���J2cJlY,l�2b�F��$�Q%R2L��dƙE%h�h�E46K(�Иe�4dƓE%)�dě�6LR��,�l�KSE����,&)��$�HdƖY,Rb�,fQ�"MLffQ)1��I��٘�E%���,�Q�bLY"K�$Ѥ��b�R�f�)"��XɍI4dز�RhH�(�Q�1�c&6H�1SJ$�Rh�l%E�E�I�ɣ$l�ĘK&�*2��)66MId��%�D�i*)L͋%KF�cJQIX�-&���*M�E$l�S&$�4�),i�	�Rh�,�4�6M�4�-&���Ib��6-%Kd�%J,�6Li1&œD�LVJ�J��,��*MIJ2TYJ2j4�6LR3bJ,�,���)�%�4Rb�F�D�(��Ц),d�2R�HIb�̣JeD�JD�&��d�IC2����!��X���Qkc�kF��"�Z6+�i*ƣTQb��lZ(�[��Q��b�V�j�m���m(��Ʊ�mQ����X�J�I���[VزF�[��5%��b�Tj#�ƬlV*��QhŢűQmF+���lj1j,[&�ƴh�E��,ZK����Z*��X��6�E��X�Ս�mb��Tj�I�6�1[cQ�ƨƢ�ZŨ��JƤ���X�Q�b�cV+I�ѵ�ب�-h�Q�j��Ʋb�ƭQ�X�*6�(ƵU�RY5�F6�d�-�bƤ�mh�ch�6-h���-�d�cůU˕��1��m�*LX�Z1��jM&�V�3E��hŢ�+�d�lQ��شl�����mQj5F-�����T�Z,V2m6�I���T�U�Q�Tͨ��ыX�lTX���cF,TX�4Q�b�ѬiJѨѩ�I�J��M�c�Ŵj��&�j�h�d�c`�J��i5�E�IE��0Qcb���j*JK&�K�,m�I���э�Y6,b�ɍ�Vf�(���ڍ��I�ZL��L�Rj���Qhыd���Œ��&J��ɱ�1X�6�LX��KF1��e*LcTX�aIF,�эL��&KI��TZfѲQFMi2j1���)5I�IccZ5Fъ(�6���KI�Ţ�EfZ),��(�2d�Q��%FJ�1�&1���س6-��FJK����1�FM���ر���U�X�1�Qlb�RcMI�E&��d٘�eh�*5��c3�-c6K�c*&mF��f1L�1�&i����mɣ��%�ͤ�1IE�Q��b�c��%�k3��ɒ�ld�j���Kd�1Q��,�&JfM��e`�LU&ɋ2S1Q��ь�&fLb�2c3F1��m&2Rd�Ō[&$��cIE�S1���Xɓh�3FS33�Li��Id�R�fd�d�XL�1�M�&KLlZ4j+%F,�Ff2Rd�6�X�c1��زF���ɣS3(�(ɓ�bƒ�5L�6M�FKb�ƙ��,l�0[�2l��L�I����*,b��lY6�L�E��l��j1�Ɋ6���4hL&6f(���LF��)K	I@$"jB$K)�jC��Q`1F�Ѩ�P!���%� M�lʃFdő,l��4a*!Qh�J#cx�\h����LP"TD�&"(F ((�J
$�l��U��A$h�RkED��E�(fŋ&%��`��j-&� b��I�ljN�\RF��)�cQL��KE���cF��1bD�Dh
6`2I���ldH+h0Q�F��6�cb#��h��1��Q�"��-�,ld��J6��BA$���RX�J���Rh(f��l!c@h�4cF�k6�`�F�P��l�,!F���QAb4F����TDX�&�A�,���Ơ�X�6+F�F# �m���+ [��BZŬcb��b64h�&ѲA`�TdōF��j���1���E���4�`�lcb�b6*bѨ(�TTQc1�(��[�Vƴm-�4Z*j-	��l��QF��ci�Q�Ţ؃lU0lV1h$�1E��VCci�b��6�ԕō"�4h���QE&�d$�6c#0�BL!(�F2�22�`�I0͔�PBL$ ��I44�HI�d1	"LJ�BF���)�	
fE3&1�c$�I(&1�I2a�LI�4$`�Q�4�d��"IID	AئA���22i!2L��$��Ȓ$L�d�H�1����"A&�	"hȔ�cd�E�#�d�c0���j&F32$����L�*L�2a4$RRh6&i�H��h�I1�& �h�S���	0̈́�ɒ�&4T���`�B2�̄��&1��b3(���{��'�� ���{~|��PQw��&��z����(�Iu�2Ϸ�r��`?<�Ǉ�B�_ {c��\M����о��ш�DU��)���_GG{�@�~��#q����{@ܽ�!�v�WZ�b�ǐ�Ϥ���,}#�Z�r����,B��A��;�gY����h���rrvX��t�n��"�'%W�t�a�[�0q��PA\�ѭ�bSa(%�`��b���G77W�1
a��K�ST�B+����%2]�F#�r����,}ƈd�F�q,9((��Cm9���>X�A� �PQg�:��pa<���}x=�CkG���XlwI�;��zG���tb�x���?�O�����=LPQcl���r� "B �R���BXO�M�K�n�9.�+�2j���\ri��v��vڎх<]��l�J|�uy�5�"ArZwV��a�s,��4up(7$$���'_�9��j���MC��!�)��9�7�!���B�Bmf�9�'2�NZϬ�[�ߨ���FGyFu����b}�8�`
+� 6��P�ꇝ�;0}F�Rm����8\(���1��r?&�D7O;����_�x� ���e5�f�.�e85�!�s�����$��G�ZeR$   -�   �                      *Ew�*�R�H�P�HT�U"�R������%EJ�%���U"$I
�T�$J)T�T�
H(����uM:�   @  �     ��Aө�U�: @  � o���QD��*�I��T��&�  )�OG��>��g��^����=�<�K��{��_{�뙦>>�In���ۛϷ{`��r��󳯾�u6�>=��������[�˯�5���i���n���j\���( =����v��ͽ�)}��7�շuVƣ;�*��`�oo��>��A���lאP������Ϩ������zO��kv�{|�ײ��p�}s���e�}�ﭾ�%0 ��  |}Q%"P�!J�R�\��
=�
��ɾ�Z���56�����z�j�������n��w�|�sĝ�ax����w�Z�c�W��]:�;���4S|`c�ov��>��f�]��P��E}�|�w��aѫ�wT�pU P� �sm޵�}��wۮ>�����<|H���
��i���4޷]:'���.�Y�o��o�^�n��}w�����Kf��}������Kd�|�z���w�a轉�ם�֗oN�B� ϊ������T�%p��Nt��]/����<{=k�=�(�n���4���|���χ�_{����}5e�w�}�Z��|m�����;���e��� +���}��v�D�}̞����|��h[X�7�O����|8����Z|�w���w�'�}J*��{�m�[�w�u���uv]�^O��/>n�϶G!���zwb7����=����f���7�����D��wC��w�s�`��퍘v�E���(�J�H���J���i��.�E����}5���H�W��}���^�y�>���9��u�����}�����R���KM�*��z��j��V��R0���}��1�z�O��].�J�}W�U[��o�=9��eR( � х����m�p=w�����<{گ��X{�+��ڝ:o��Jk�=����<�&���r��I�C��}ǟ`}���À @���%@��
"��  �N(M��_v��j绷����z�շ�x����=�R��O����w�X�r�����{��������s�Y�����|��v��8 
 ���*O�z�ǠD����+<����w�>����v{��=b�\_@����b�5��T7��Wy�׫/_C<��w z9�^ԀX��        ��     �  �� �J�Ҁh�Q�@i� �� ��!)*�       z5R&*�OQ�`     i�T�
�P�h�  	��JzD	*�       �*��#05 d�@�14yO��ҏ�~g�?Zҟ�Ǖ�@��� ��%�V�� 	/��(�ZI	�H@!%LI����I$	+���{���?������t��W���>G����_`!���=�l�IJ��I$�@��C�0�h��?OꁦO��P~,\� |z$�$��O�?����/�����ؐ�HU����5����/�[`~�����R�)KJP�^���y�BW);�JeQrq��	?H$���w�[����Z�	yz�;ަb
�o�#M�p��Ӛ����.���(�fp��(�no��r���srYn�.��x�5e��M��fP�> �>%<ȑ�2�\�M���m�I\i���t{��J�"P��m�Ge�v��Z棭:˘���t�5��S� S�<Mr�@iTR�J�)����֞WZ�����o*C	��\�"�?��M}8�$���z��J
�\��2\�#Hk�����*4+.�����B�� �H'��޲0�hkU�.�C�`���r���:��G�c9}OԒO��W>��vmA]��o<�	zz��9��OvCmN�d��]%-ڼ�6��i)i)��9��˽/7p�Z;!�:�D��K���)*|h�L�4��]kX�k��a��w'�PF<'�����+�'K?}����_g��8��1��q�����7�c���=H[���zi8�#�P�P�\�9�&��w5�mV��/r_\!��!�A��1&��Oj݌m����)�:X����IB�qvc�H�1]T�_}�o*4J�;�4�	�`]�vb�q�^�zE�l�鴞�n����T��B#���i:8fF�:.��Wr ��Ը�����jS����qa��/�>�aFH�?���3�7�8.��-�^�!? �$���s�*� �ךNf��tơ�3{�%;�iCM���9��mq\��C���d��cǫ��ۺxL��>:�W9un�rd=����[y�9���
!I�n���H��D��sA���N���+*�R�Ÿ��"ls�,�s���'�mS�	�E�������Wv�LM�A�2�H!�4J�qfM��e��fRՀ���N����xܧ\�7g��R5v�ۭ���x]ᣣ]�1٥h�dF��%s�?E��Fg=�ƥ�$��$Ou��d���+�]�I�t��Y3�!Ճ G�N&�q�^�N-�đ�\�g!"wR�W�:
�$ɝ�Hçָᘞ���L��L��~0�흙dqQb7�Z�B�pʑ>�)?���ե�a)5�*%nq:���r(LolO1d�#���tu�ۼbo
�Lk���c����K���ζ)���D@Uě��[r�fr��u��Ǔr.$c���!�9��`M�u��V����&��+����9n�Aޟck�K�!��뚎���z���l}���g*Ճf%�>\��j�ę�\=�spcI)$�q�Փ�ALj�ol�8��f�*+�� �{���L�o]�|�&��ŏ4E�r�5T)�gœ
�J�­&���#�:S��v�3���ad"8��!C�`:���	ʩ��'�?k�U�Sz>���:�\^-#w1�0z-��EЉ���r���l��<7�3�2j�/��mE��V�:X!�+��h��i��z����K{,�z��(������v�-����iS��JX'*F���aE�����/jq��D5=�6u�Ou2wr����_�H8��J�q.`���g&�b���p#*�P�eJCsm�Qg������&�����ϥ���C��&��53��]����� 8���R��K0��zvEpe�R���#�.���[���zS�i�\s���Gb�bIb��5k�H,M1�]7�[�m�,���w�+6-=���_k�p!Z��q�x�Mcye�f���2i���BY�����D�*wPh:�VW2u��m��H�Օ�ɳ'}�I�,�GX��-qMS�ƳtI�������.q\�h�,n3e7�e��K$��I�]F��R�bF�[�s70��(�tR.���nc˙����Z�fHX)�I'Y��i�г��6{t>2�c�l.��5�2��f�z��f�)z��{�f�eк�sP���bT�b��f-!����c�r�7n�9���i��,��-ec��2)<6�~з7���M�8�8�hN��E�
!4�6Q��.B=���ǹ�k��7�{'j�'u���P��L��+��5��;��ٝ��������ܺd@�'L�y�i\A�z�F��P�E6��,ZF�����Xې[��	 {8��Q;�=AK�N�vj�t��[�ڳ/r���v�uN@�n4n�ç"Zy�i����~}�%��c�j˒�o���L�%�dyaj��լ�_`�ac3	u�?���Xq�Q�3�t�� �fK^�ǽ�éw8��ro}v�M��'z)9�{Ǟ,1��sx�X�{�gn;�sN""�m�J�E�P��˝��8nUv�%��:��\+\�l{��/	�Y;,ղ�:���]����6��$"�;��2����%�;��>�!�o͊z�iK��r�#:��%}�7�3\},c:�w��,��6q.!ԝ�{)����V�f�,|�kF<pF��t����q��T�P����Fv���&��~�_}��j�Ys7���3�u�o<T�j���>4����w��b�����].�tJ��#tpd���w���֘����Ŏmt4����z�q�T�̝H��;p�l�F�܍���Ⱡ��;�Jm߰lR�J8��T���&̏2<�n�=���&�˪����əz@������i�S� t��p��?�Z.�)G^���� �~P�~�Z��G���s�r�����$ẇ̓�<��[��r˵|H݂<@���[p�!�.<0��Ⱥ����a��}t���������r<At�P������)���Zr�g�fb��·L�,�Y=2��~zq��Z�7�9P'�GjB@�4	��?3�9cDS�s��hS���H�;I5=8�{Mٛ8��w�kHmG�쾽�UD��dL��z�W/$㗢Qۙ�F���֬���V\�7W��1VIJ�i�6����-���3�k!�M��b2�v��JuH���f��Q�KB�Ef7b�
��JF�GL���ZQCI�����a�H�i���9F�-���Z�$TQXgd��O$���ħRF�ˇR{[�8��Pg��Τ)A,f�Uͯ
,،[�9tMfu貤i�`:E��Z��#�SƖx��Ϗ{�!���NSܣGTi$��T~|�=
��h��D�8�-�m��>�'Q�bz����1Z��=C��t�w�<z'��a�5=[�U�tC����P�b�����&V��_'�J*�Q�j<�՚�\Q�=�*X����F���u*�]�ya��i�B�t$KI}�b ���g+�\�.�)`Ȉ1WŴ��
jP�p�Z�P���%&�79�MI�H��"G5jꖩP��⍋j\�<y���y�%��Zzk(4RV������^��/��Al<�9U�ĹV��#�qF4��$�$�aS:N.�r⼺'Qk���J�*�jڙ�lt�i�]3V�yE��F�Ɯ��E�3�T�q����@p�e��F�yr��}ʹ4�oK�gf�;y�����q����$�r���R؉Õs]��ĪOU�j�M�*i<@���b ��Ŝ���i�jò9�CK�*����&����t�>N�DL�QC��$,U#��x���df]k�#q�\nbd�K�MH�5��K��t�y�K�J�p��mv(��ϡ�lx������n'�I/��R֍Yb�8�U/�5H@�SO(�ռ�$jj�5�{�ujR&�kAmq�qv����BvMEt��sQ�u5�,�4���b�E�I�į[���Mh��t^�t�ݫ�ۋ3.��.%�4���"t����N"5ذ�9�L��$I�[�W�5�t�Kؠ�F1w^�����qK��؜��jN<;U4� �H=U�shL3�#6K�Ir-���@�r��E��E�Q,ZFa�j�&���M���m�6��#�5tIY���d.�B�j��xc\�ӅiZ
i�ƥ��]a��r���*�QG.6�Ӊ*�fqmŁ�^�HdL��w��z{�{T#��~I:��b����ċ=E��,�Ī%Z����!��R���P�&���h<�o�]���ڹ�qn��t����n$�ɬkߺ�'Osv�s"U��B�ֵW����r��"=��ǣ&cb�;[�T�[mģ�1E��F��rN�;9���ͳn�ա�c0(�&�c0��<��9:�o ̩�p�0�"5uor�N�ܒN���j-Xp�O���?i�~��b	sک.0�(��͌����lc�n.�죊���eN���Ovq�t������.ؚ)�Ƴ�t���kA���Y�Uq���D�8��5�qx�E���\to>����έ]sv>V��6b��՘�O*�/b(���䁐,��b�5�Z3�{�]���|5r�\a�e��]6�{����H̯C�[��#J�3�Dy�o�oW��jڨ׃gvGx�TP�	�on${LQ�}0nn��L��{`q�͎�e�%O*�]��Q$��Ž66�ͼ7�$:$�k盖�&(�gfa(H��k���U]D��b.>�Ӄcúx�	ɧt���6ٳ��b�N$[�(��kc/MhX�}�f=�&���hOr�6vcPj�h�$n�jGAY]L4(@���dUb�^
���ƭH�G=�&50�����d�Zy�rg1��u�َr��wzk�n�Ã�W�:#\mOZ�;�|z��X��m�'%:�eM�\�p��u�Æ��M-������;Y������Q�y�ېNV�s�۹��0�#7�G�p�ח!�U.b��Tn�B��ㇵ�6���L�lě<%�n:/(���kH�2kP��h1ݥw@�xN��<��V��B޽��糠'���429�(�7{h3���O�ƫo"���#oM�o20�.�!��Iʚ��@g`h�2k�"{�Q�1����3�Z�=;�h��.k��.�g��wqf�v�ٶq��s�K�<֧}B��y���M��ӯ7��q}�',�n��o��1�dBw��gܲ�:&֧�A�C8Q�*)�W5�Yθ��wB	!yQ�7�N�o:���պs�u͌k:�r*,�ŕ�5��N�bU����bc����a�o9m�:N�_Q��E1a\{3�跺^�S�%�2pr�$᯴�fu�Sjp,��u��%���8#n�ZCb[�JX�ᝒ̷��=j�%��<}�ٵ�.�#/L��%��p�"���g���J�o@��Ǆ�S�3�dR��\��I�Uvv�.kh����۝`�.�5߶f�C�f�]���ާ6ݚ�1��f�igu};ff�
cz�(p����޷4��쏞Õ34۳s�a�J\][0֤�50�T���s���Zy�s^�t�e��cI��0��OM)c�)�uX� �u+�^�]�Zn��G9<�~8�Ʒ(�Xւ2'ݮ���:��h����H<bH�4��Us��dUv
�N�^:I�9�K�"P̯~�Pz�Ll8s0���h&�̞Ňzc��N��ר��sJṚ�c*-�I��i����q"�s�v� �Jw�c�.�[x�ץ�¶b�-]w,��S�v��ơ4^j�z��(���$3����3V��J*u=A�.׋����wvG/}G(���-Y[Zm���;l�ö�V�C�!))w��v���`���r��"�Ȕ�V>�ɣx�},Nf��ns��>��c�2�;�xEf�_sXHy���7HF޼��/���!44˳��̯�4�����j'"U�m�`B���E2;�(꽃nq��I�x�s&1n���N#ǘ$�6�y`Θ�Mŏm����]�Vt}���,1�-ǧ,�S(Vby���5��GG��M=�D�k8�Ԗj�M汖�u�=�=�89�3_QP��tv�6��4˺K;�t����3���o�,�,L�M�1�$���pVL�f�|�E#+S�î�r��={aK�{fn�}�c&�h�G�:Mᓤ���oy��{�`�ݚĲ����v�k$ɺE�ɑ��D�fdDE���-�Cٙ���Ŏ�^+���̆��,�u�C��u=X;��L��ӻ��Xo6t�i�#:�^�c�
JzD�\��.�Q̸3֖�i\�a#��iؕ_��êbkh�Џv;����ZT�˂f>X7�Ֆ�un^n�5���ns��+H��K�S��	 �ծ����/�m9Ǩnq���LJ:���z7����j�hPUQN&:���EZ�Mi�F)IqF�V����:�j���6���̐�cǤ�2����ι�/�Ay�8��u���Q��n�6�Y�&�T����i�Z�w.j����Ih�yل���'��o�a_��_w�~}D7���� "�^�� /� �5��&D
֘nZSWl�h-A3�2�,ع�)�,\��t%�0�:�뉦�P[��ܹ3M�V\���]0-�d��!��شk�1���`]-/h2Z�ݔ��a[b���Lʥ�Ц���t"<M,Wm�Y����`��R(b�dQ04j��b'R� ٳP �kf)@�Q�1�k��ĪJM�8��ǒ.�Z�c�s-�An�iM���P���ua�[��ܖ6\(7��{e�0�V3(�J��K)F�z�uL�7b7CHMZ�j=u1rk궔���v�eu�/�a���f�)���
����0�@f�wk���#f��H0�d�3��k49�{/c&�4���R:ڐ��B�R1���Қ7K���R�Zg4ql�R�[r���Hk�H���J��:	Q��Ȍ�	�W"_(�Yt�X#h��Z�c�c��4�!��ljVe1YiB��ka%�@F��m���C[���m71hM7\�Cq0s�J�jA6�@�1�IHY���D�mf.�!0�,qST��3k���\�Wks+@#�T�t���1�^]mVa��ˆ��mL�ël\ظ�`xY��i*3r9�`�0�C�w &@1��vb�fu�^�K%(�GT�A�JR�F.���k0��m5�I�𴧉44F%ttW0]V�:��#V���)u���+��n�]`��v�tő�Ԋg	�Z�c�bV��j�<��f�ҺP.��֥J��n�,pQSYlrUK��r��.�Z6���f�`�K����@��k��9\-&#ΧC���Ul�2�e�-e�T1�޲�R��3oj �Ê�;�x�1���i��J4у�ҕ�f�95�����e�,t.��^ô�+0��y�69¸M�&t!�5�jg��J\\YP����c�kjJmZ�\T�<�����M�Jb]�]L�rq34�]�uhl�β�\�+aZssk��k[�a��:(�FT5	v��+q4�lH��k
�5]�\;E�l��p�`�sb���#5��G92�a�Cs-�l�SQ����� �M�f�Jml�+e3�ˬ��%���3
�ץ"�1�Z9�3�l� ��3;Y+�2♚��"���JQ���W1�s2��K�Ni6I�m\�cbY��p�s��;hx��U�������%�ŷR��ي���]�Y��-"�DL�K�����P+�L�tͣ%�]�0����%dxb.����b^6�u��)I��X�e.�u��P���GciD��c3[6 vZ�	����L ܭ�H[k&֙K��1ř[�9�bJ�80D�/Ke���4-[�Zj@.�sK����v����-a��emcІ�3��녥Km�_<��ɍe�E�J���B�F�,��D��.h��FZ���)s45��`�b�VҲ��!����!SL
8�ѩ$��aƺ��g9�iTZ�P�Bj�JUḲ��\��2�c�݂�#��5�`e�q1V�[V�c4
X�Q@%�&��iqC-53��%j4IH8�W�[	�]W-%]�nV��H`�#hdL��Y\��VݢF�W`3ăй�M��(�sY�l6R��v�؋kkM5P�r��n�n���^+̡�t�G��ܺ#rܻ�A�����8��M4�ʀ�**��E�:<�Z�m�xF�+qn�Bܻh2�aX�k[�-c[W&@#X�]0),s]�3��ѵ�&����&Ǝ�˵)�ITeKi����c��1$%�Z�0M[B��&\�Y0�ͮ�[r�\�Z�u�Ґ�-%��%���B��)a  �em�ղ�4l�n�k�]�n��.�a����3�-�����������h]0�����孫Z��M�tX�2G9�ۄĮhJV2�JV]1^��і�%��� T�U1���b�.��6el���t,��5#.�W9ݘ��:8�mr����'���J�z��j�&x�� �[s-��)mLԚ���FL��:%�����][��ՙ�0ܴvn��$q5��tXYhі�e�%X�u���a�m�Ԕԛ�����ab���v�m����"�4�*�c�ÃgP �L�v��ݨU暭%��"�6��&b,�f��l��M7X&Y�u�SM(�R��T����cn
��W�����GK�A�w[a���n�����-��[������[�7����MJGQ6�� ��SAE�s+m!��ٍ
��΄�a,qz�QEf�X��v)1���X�&`X�����m5����J1`5�Ƅ�&4HF���L�,����&1qe������:�e�XF;�ˣ��`�If��n�q�fP�:mG�\l�䖠"�%�8�ƈ�-I+2���S�k�L#��a�cJ�XhEَ����M���e�h�GR]���:�-��b�e�le�i����ֻ��/��ګ4WX�Ld,]x�*E��舫M�tCX�<�㳦*�ΰ븶��e��5���V+u��5I(:jd�4�$S��F쒛X��*&ku���Ƹn��%|/�t�"RGcL�U;\�\�Xb�Wf��6�QnjY�%�FW9��iRUz�3�a��j+��:�Q��#�����-��I���Ք[�5A���Ǝ�U����[MJit�fF�V�B�/�����[������,AĹ�=l�V�l!�#��S^Ŭe�p-�e:�J�L�k���V�(�T��b��q�]��6��4!V`lI1b�]iF0�r�m�,��X��H�F�pV���)-�&e�cvq�PKx#l�&
�TYR�h��f�BB'Xb�Ʃ����K%ˈ�up�
��j�ع�cX���m��H�L$
�F��5��d�E���j��b���O!1l<n"S`aq�mMu�+���m��,�0��B�.H1hu-��Q�XV��-bYs� ɺ�2f]3�e��YC9FRJ��Y�����y�v����qrb̘�7(;#DqͯV6��+�z���X�-����+��-VnQ���[jBg�#�&u��f�ՍqFZ@�����a��"ض�HX�9��@���ZI��Tu�K��կ:=�L�����F\%��+�1y��V��SV�U�f��a���ٴj�*8�t6�qCnĐ-r�R���K@�S�K�]���*�tט��*�ˮnZL4ИK� ��P���2���6fm�-�����9I�XU�X�#e͔�6�\��KpVYu�"1�٥�L�@�����h���x	�^����jb]l`��̋�H٩����A핲�Y�穩!�����b�31�R�7LG� 4�چ�M��l�o]sH���B�U�a.w��y��5�4�^��k�� �Y����"�V�V����dƌ-ؤ&�.n+G"46�&����V�-��� YV,"Xؔ�cA�]���P�oXG8���m��rY���qs�!�<^��1�q^�F��Ak+vڙ�����E ꁄ�-��!���]/li���lƁl豨1 ʫ���Ɔ۰�me�ه�F蕱�m �l�%b��̸{S��rbՆ��9��gF	K��L��)`����e�M�P�ѭQ��C*��e3��e�X@A����Ku�Lʹe-�Gn�]�,-�*B�R�8%�6@cf�j �����i�6f�Bꅮy \[��Lױ���K��n��\�Tp�X8MF$�-[y,G]a6��m��eKI�F���RM
A��CV���.�n��&M�M�VQ&ғ2�@+7YQ+�d�k��k�ve�a�g�Wl��1���Yt���d(��:��Y����ch�)˭���bڳ-lщ5�,t�$�,��3^)��W�xb�`��� ���f��@�K0�Zk���%αv@�6ԙҭ��q�Bk�j9u"Xf�\�JKe�A�U���k�y�x�:���.Q��X�(@�۵49�1θ����6��t oYD��Q(KU��6�&���)�3kV�9��l�C*Gj�9]H�������i��eZ��KH�an�3��4jFbF��q1�e0�GTG`�t���^*9���]am)�+��)���\�+�u݄K��a3f�dux�%@�\5Ô��Z.F�]o+KQ��:�J"R&�910q�17!�a�X2���Bl� ݵ��mb���@#v�bI�SJ̩F\�����Z�4�칍�uT&,��u{��D�X��&�m��� fP2��.n�(&�+,3�Sy"Q�ؚ)6��������\��b(�B뙍x�"�f5�
�6�3(�kN\G=vlt��jo��F�y�q��4cV�K[���v�������١��C:YliR�.�)^1�)��
����-���<�,L76��Sia��ZƖ�+eԆ��A�!aNjbҨ��mQ��k�b&L� ��Pe�ؕ]����5y�f����̧VW/Pй�#�ɫT��R iPI�!X�&n�X�uئ�Q��QKv2a�"�q�em����&�]V3M�VZ�2I���ڥ��)��4�B3#��.`&�+&&,@�@et-�5�&QQLV�.J�4e����Ġ�@�֦�ŕЎ�:@c4֑*� ��
P�ض0�Y��,^ڻ����<P��с�CifvH��l�뙰��&�*�Pe,p�-A��R�]|�mm:�l�V�܆+�6�u����:E�A�P�jں��0���3v�˖����aٌ.m��mJn�U�ԁqT&,��.Y�K[�4�g")e�F��fk7nd͆��3k��:ƹ�3 T����b*�].n`�`7*ń��h��Q��`-	���q4fuJN+u���ɐ!̦h@��uT�2��ɠ�b��61��Զ0��j�h�)a��]M�f���3���Itڴ�4��76�lL�EF+h��f�W�t��UW�%mΉ2W7$ѻGV馭Z�fĊ�-�v�
�F!�.��{J��܊跌^a6i�F��[���+� �$�����Z	.���k�^ �~��� @�/��g��H���H������ G�b�򀕴��zi�b-�Q��~{�č��TK�H�B��5��m�F%�O������֖��B�h���zk��?�چ�H늙~�L���j��#�"�G�Ɵ�y*/p��2	1��eP5wUɒ��W���#%��J'󺲔/�V�*B;=C��x��X�!����H?�_D\��A��k.�@��7�=�/iY9R�s���s��%����~�߇Zs����eYׄ�b�S��4��x�E,�UzwCF�%������T���~���-d� t�w7z�{7�8�H{�����Fm'
�^�{ �w7oP�B��i����f�sU�>S��pN�.Tl�qP�����Hx��V�9����Kr}�ۏ�/.>�>�Ï����R��q	��1�c�Ƿ��'�=w�����a��p �1V=��C�>c��2�,����Z5����-��S�_-4�� K�X>1.k�w��Og��3���9ɼ�`Wc�ų���b�xW�6X �%�������~>�|Sv��s/��j�Z��X,�D��vsi���ĉ;;��5�sX#�K�hkf����r���7��~0��~	jb,����0���O����`]�ݺf��_��o���(|.����l��e���~
n��J�؟ؔY��.j�|	B��g�%�4�����L�|����0���T�����2h��u
�h���pϦt�9w����L|��%���,֪�|8T��L+<�>�ϭp��=3�n��K���a��h�;�B�^��z��x�kA��U^r��p��B}�;3��T���������o~��Y�߇=��"��b�=>�Z��e�Ì��f��r߅^!0��\{�M�=�Rs7���>@�%+��r �L�&�,̂r�Eϱ�͔}ٝ1�����r򰎶�.�=��{)�wz�6ɾ>߁^�ve��=�:|3�~�"�3ʵ��"qy��n��x��a<��{�"=�Z+X�0o{�L�w�^�!���'h;�Ꟙ�l9wN�n�����9>������?ৗyAbOٷ�?'�>7���v�	r+��`�n[��'(�&n�޺¹��'�)��o]��Tb�x�lZ��|�������:��r���ޝ����1>^O=�i����^q�� ��\.yBe?d?1so-���@��8f�]��`��Y��9�f���,�ᛅ6#��^enS��(G������&����w�Qj{F?�R1p[�;p�~�_	���cG���p7�bG"�؂�.*,��'ƀ{�dD�j!d����{%�Wb�R�꛲l��7Ҷ���=bŦ�����>m����v����J_5��{������<�>�vw�>)0_`���	 �lG_�vEGڳ}<^�yO5����<�}�g�S����>WM�~]�(<�=�����q�`�א�A���h7�P$�`�<���N��I��Ϲ��Q}^���/O�1�@��D��Z�6�p�9�N|�C�T���}���nZ��ݾ��X�2ź�ޛ���M���.��>��>��ɟ_n��Y�����\��=����
��V�.£k�fb�����y�
A_� ��o�~���~�`�Z�x{�{߀L����Vf��_��Y�����>��'�6ꄩ>�90�κ���>�m��ʖ]3��P�2��v�����Ҭ��}�z���B�`��`k�.}��C9�{.��\��M�����q����~���ћ�8��G�*}7�Atm���M;�EB0r�Ј��42q�O�K����8��N���ݽ����nu�0����@��ӵ���`�4��H�J[�ndÀ?��8��I�-�=��(/8P=��n��7��~d9���j���J�krz����o�E�J+�x�6��O���H��(2M�F�'�L�cs����'���Ln�Y�>����w��s���O�B��Ȼd�r{��.����sy�Y`wh��U�y�AN�2����~�m�;����8,��-3,�0c��lX���s*��TN�F�\}rY娻��y�zm�_@�GHh��/��w��{��Ϡ��!��:�=���/�Z�5f��� ����l�_{Vn�S��`5<�߯�r�f����CFhDOB %���
��u��*x����T}�%(�"{^�Z������6��&�-$�L1��NK��wx;�I���}������գ>�Ph�!��K�|��D1=��|}eK�Irw�("�ɭ�b)&�4M��ښ�.����0��n����@9wa�=��}���tA�^�w��'l��/���۟}\'�3��=�~�%p������эOe��
�e�<�r:�F��u>�ȝ�/�`��>tw���~#y���'��a�����_��Y�T����x7��|E��_b:���xm̚���^����X��t7ג<Ȼ���<=G��Aˈ��DX�-0�o9�֡x���K *oޏ�/u�V�w�^��0_v�u�<���(ݾ����o��ш��;��?��$����ߌ&n`ϳ6���1�;Z@L�(�c�������DD8���:7�-��7$�h��v�=�u������,0��H�Í݆�wޞ���C��>����1�=���>.�Z����H�}�M�� ah��'�a~Cv���9� ��~�T��Xn�{�:`/�3�Y���h�Ȣ;�w��|d��g��GP�\f����<�E��Ės�7����>�̃On���F9��`���[!:���3�ig�I�0�� &�F���r�X���Usw����}�t�u+~�m�{��s'���l�ϼt��:�sp׃tN>���=K~���n_�����ϲv��q2��n��ɽ�hX��I���Cރ| ���@���`}�P�]3>���>:��6G��ﯔ����A���0��>z�f1�\���,�� h�G�J�3��+�d��A����W�>WW/�}]T1������ݛ;ۛi��py���r�χ�C 7�a��9ܙ��:{�����M�����:3���C �<�\19���A���-��<ގ�K���cK��y�Ico~�l<��z� ��w~ˋ�~�X���"�,�ev���ۋ<o�d�=/�J\qϾp�8 4{����>���zw� $6_r�=Ŕ3�=π󈟵&�{2�LK�� aH�S0?�>�s>�?tjg�(�oT_;��ve��s�T<m�Q�yol��c<��P�g/� �l ��΀6���7��.���� ��ܚmaI�&s���x"빾e�n�����ń�H>nf��=�3�.�G{4�̫�!`�޲�,�맾�����o$�+�#���=ΚpK��S��G�j�=��=�|�j^�b��cx
��J���t��-_|7΃g��<���=}��.CX���t�ڭkxbF�Se�KO��k@��_]g��@}y���� �ަ�v�6�ys���T+V�Gsy�|C/�H�
8�� %��3y����sy�ٱd�SUɼB�^�KV�SZ��л�����bq$d�j�P�f�Y�6r��7�현^���#��ڜ�@���.���_�2�TN�Լ*��}�yE�
�H=�+�7z����� �/,H��r����N�%��|v�z@���7�`
(�+..��Ҟ� ll�6ʚ�����@����_8�`+9���%�����æU�HE�ޯ�I^7n��w4 ��ޚV�+:���9��|:��HA�G2���x.n_ff�� �r�k5��S�k�@fd����A�39�A\�%��۾��.�ݔgNN�\��Nh��BZ�6f�Z���#�|�#M��i#�Ν�o6!c�ޥ	��֊B2U���jl��_dHZ�r�E��<x��2����R�m� e=��Ğ�;bZ��"�s�Ѫ�������@�S�Y�TT�H;��`�I��$_9B[덊����r��o�#g8q�o�^G����>'h�׹��Rr|9�x@+�����R�M�����w>�6<$��肞ռ���Y�g;�7�c2o۹��X�S�y_�Ź�����YC��y��xgOHׯ��I�w�����a卵��xΌ���}��B�_2`�����Gv8z����ڻV�fL#7���;���ΞWx;^խ�p���ێJs|�ً�e�8��]���N��n�y�Y�/�O]ZȺ�\�xzZ�rG�3�n��W`�?I.����`rY��xP�-��sϻ|Hlyd~�7�̕�����=(�;�#�<�>/�l��s�Og̿4���Ӑ��L���De����yv����m��ִ^9��y���M����;�aɏs�<�V�g f����m��Co4�Z*���\��������ʻk�1	�M5^�Q�`v�j�]v1�s�j9��	/��reɞKy�/M���->"�/�tx��e�:�é���}�;�(!%��Z��GYIw���H�S�J�ΙIGs��~�׫��3�P�?K��07��s�Z�}���'`��ݝ1T���%���ze֊�.�k����
f>�4覌� �[�;�t���زzC���6-8\��ޛ�h�����Ƕ��1J����(&QXna�q�.P�x��	+ZgD�t`�Î�X:mU~ע�A�0��@�}\%��>!o�u`Y����$�qSv��/qK��<�`�w�(��HG$S�*h�{ٻѭ5(��m����\ݝ&�k��u�m�z}�������e{������a�Gj�w_l%T&U--��}��q��g՝��.����4�}��jY��"�#�}��&Ѱ�0a;�d����?\͘�M�G�<.Ỿrw0�ɞ���g�3��_=��E�F�=Ǹ��.Q��:��}��'����|�����ܜ��	�p��̻h�k����9{��z��k��������R���a�n#����HII��-�/��aC9����3x눙rWf
�څ�e(MaE�
���Ҝ�`�L�L��6�y� -�!Xs�h\8/f,f�
TR�h93m�����X"Av�f�Vba4�x�RV��4Q�Jb%2e��1*9��)ut��r���t�QM{U���M
��[U,v�7b܅	R�5a�4��Kw��̰(��L=��.�l�A�8լѳ*g)u�نc��3�]2*����[�ɕ+t���ة�����]�4�v��c��+.)�)�,xI�cS'm5֘�e7eԹT���BJRZ�X]�X[.s�����:���dC6�$��5fW;#��	�ZMcn����ӝ6HZ/iiD-�u��G�c4ɖ�"���)-:ġ`$Uh�u;Ե�/���e���&�u��m��hŵ�e���L�I����&�-��"C�A����j�9ّ��2Ҍ�c�I���F�Z�4��X���!�Ǵ��+� ͘�.֡B�]NU�ˡe(�Xeu��k�[�ŖV�l@![��e^��d�#3���l�e����q������pVX�4lEu	�%���,p.�fᄢ�u��-bY�wT����6	u1��g#A]s-�4��]BݡYI�K���lƯd���m�f4L��\�6pYI�MpcL.؈�P  �(�\��� �W���قB-�5b�����*GZJ��5����j�:��;6l�X�Y͢;K5�M�KIhl����ɛ4���a��[���:��t9��EZ٥�/]��[�X1�]|v��<F�-�I�`,6ˈj�Ըõ.��F�HQ���5����"��z�����Ŕ	m�.)��ل����vVl��P�#:�в��V3P��Fh�C/[m�E��2��b�k#�HUR���M��3e�HBS#0�G2��i��\!G�bJmi�f��ļWXb�)��c9Մ[:��	m5���/0�	J��*SM�]u��2�$���n��{:t��	%��4	S�*�����q)Q&��6���lK���C cHlhH�	�V1bK� It ��# lI6�m$
�v ��m*b%D���QQ�U�����Aָ�i��i���U��U��T��D�ACmQ4�j��i�r�\�bhm�\��h����%�ݩB�B�v@(�J���4٦�b4�u���2�%ģhW�Z1
1�F�*q����`[H���5�-_i+g]h�Ti7*�T����y�pJ�Djrj��Z�'��o"X�h��k��o��[@D��UlB&б�c9q*hV�b1��mSA��ASL@:�F�h[hE1i�D�Th!DA~E*4UB%q)Fi.l�"�F��KR�ib ��[HD`i��$h���Q�' ��Ƅ�� �HJ1`��� :�${�$c�m����%��4��I&����E$�rTА�q���i H�HƄ1���LH�	b��F�!�F�Am
�F�M
�HZh#IjU(���0[{*vV��VN���z�]�}x;}r�m8����Z_e�dw�ֵ�y��UV�sYb�iltelv3���h�Ƭ(�b9i�9�v,3������ˀ�0��+vR��M�!F�������]Y���]�p`Բ��lJ$���`�%uņQ��ю�&�S4@3,�EN����;b�r�5�e�1�h\�ɦ�]n�3�Į��K�6YJD��8LҔ�U�(�\��--��!�l�jڮ&JZB(o?����{�N�'���E�B`�h�F�P���qy���ZbE�K$���7�ڠ
P�*�)bS}s�X [��؄.�}�hA�6��i&č��^� �C>��"�*"%"-**��*҂�

(�"P�)JR҂��AQQUJ���TTj�TDE��a�4"(R��"�K@�JҢ�%���j�Z�*4��B)H�-*�-R4(*д)��1u�e�&9l���-"(*#�%R�6�F��@�cB���EFB�ڽ��tҞҩJ�Z-H#�ں�R�Ai�DF�T:�EF�/>��ƍ��-
P��c��Z�Qk��QQ��Jj��Ph���C�=tc�Qk�D)P�P)B+B���)��Y�x�2e̼�#��AC�"�*(��騭�3_z\��KB��r}u젏����׉��Cu����Z̫��"RЫz��!܃KJ()�h��[Z�JUQN2��<���̓d��`���'�;�:�*4�8��Zt��j��nN޴ӌ�P��������_%sr+B�c�a�f7�C�����GF�4�{lk���jW2�����=�o.�l��,�tm6+�P>�h�k͖D�8����HІ7.�h�/`�IiE4Əw��{E~xj�+��W��Xqh4�J,:�v2�����T)UTZ�P3>3k.��0\�b��[.Bd�1��x�8f�YW:]�i�.�4cHX˵�V����{��;���Z�7>uj-x�Q��+xKȵ��{���9H��h�=]��^N����ű���3;��:֞��e^3��r�ܫ�uV�-���:ֳ٩��泶_����:\N&g��S:��6p=�w��\"G����D�-��)��Z�5Vح��������z��q�UI!Q{�ί@u��Yƺ��B�?u��q\��\��5U�R�̤��}�6��"��ZCsz�ؓib,\7n�b�����U-�bV�q���Z��$Fu���<�ٔ��t�����w���c�:,U��lƭ��}�s'P��jo��U��n)s�����+�R4s���ZߞZaZTS�/�0���u�n^�ѩ�з��D�_�m�oX����=O�u���|�k�]�8���s\sI�9g��+m�߯� m��7e)QK��	q5�V��u�''\�H�ҞԷ�K'z֚h`4��s�OI�����&�Qi�r���Bh�T���
lۮ5�uLWK�͢�cYtRiX�+VO��i]H�|ӿ�MW���+b|���:��/΋w�o<�F5���u�K�H��'���٢�/&dȲL���43l�3��=���׆H����y�"�"=��30^�hL�o	fK6�?a_��\���T�2�-(���;�H��
#�P�ľj�c\9������/����ܸ�8�����d��qZF�+V*�ùaL�K�:A�:���DZD�-�ĥ+$JQ������Ҷ#B�5Z�M>Og6�x�,k]�l�?e�38BS�����T�٨�.��t�����Ou'O>��˹��.���@[Bm)����`���֢4$	2�ڜ��bA���"�>�z�����&տq�����\T��Zj�>~}�M�M[����Di���o*���2���cS{�Ő���~	.��7�厯Ҍ���nҍ����1�+ve�������6��x���2%e��Xf��*��m}��/��ǆ��5z���!W��D��dq
	�M�/^`JI��V��C� �ZD��$�OD�}_�J:Ҿ���� �/H�����#�8@�Lv���m-��l�i��.�j��I���g\��fH˅
= ����ښ[Cz"B>�f������`d�,�J���e�=�>k�5t���eHI�lG#FD`H(���9I~~���+uRG�9>q<���4[ ������!�
c�����0�~�eq�;�v/œ��"w`�'��`،d�)^>$@k�",�h�Uˍ(�TH�軝d'y|�u�����B�8UR	p~A߁�=f{��'���}��W\V�qqM�^(07l4�v/]�C���PQQ�Q�)E
޵rz�\m5�H5BU(��kؿ�V�y������t��:J��h.}�˖(��avmX�Fgk�X$m�G�k64q,"u�	���jٜ�֙df�r��_��$�����&�C��J��W���_��0n@�^Гk����	���d����n�H��א��̍�'sˆ��me`� ט��sq�|�4�?2�=|k���Ë:�`qi4���)O�%�"P�ɧ�9~k��E��>bN7&L�c��П�����$T�Ȁ�8;���P{m����E6��^.��%gy3�\��[P�x�;�T�{��f�d�x���ns�2I��궰�J'�D���G���H�����"�kկ{<h��^?gK)�P���M��N�ẚSDP`��q���7�5���s�@���UjG��a�>x��\aq!�mf2Xl����V�N�5��^�\�ۡ4��g!�K)�8�L�CL36�q�6��%K=��WCt�F�J��[�w5SX�.,��,�H�e�Cc���`��Kʂ��ak����%��t{$a��&��Z�\�V����ŷU"5LQ��Z֙#,L�F�GJ��t%4�i�wmi�ۈg0-̧9	��3QV166�A+0��³E���R���lt�kls�����qF�@�F�X(�_E��`�������C�ș�;M��m3�f�pK����	��6[r�T�hX:`�{�'�N����ޖPQxɰ���wU�3%��F�Z��1�`؆4��A�u����Vi�wb���8.���ًU!,ԋ���U'0"��(@��a-	��~7��<����]�A���x�ii��"��{6�.˪�$���aMA�y��{���_b\`ĺ��ٟ]|�q���6J�����^3����x`���Hd��Mwz5�D���0���=�~���֟q��F���^�[I��B�X^К��O�D`�د��SO�e8�t��ʳkn��U�I��af��iq���`�X1)�h#{��p��rp!���|Jf�� 5�RP�t�)>�.`��\�s�X��[]	i�J5h۬2Fl7f��0� b;60l�u���J�;��2��wS!3��� ����9#ȣY�u��O�=��=�/ь�ķ�@�a�Jh�v���L=�,��+C��)��C��w��B����@��� l`�<���H�[�[��0�1�>b-�ll�HG��G�y��i�B�$[Q�y�o�M�����K��3�b	�ؕwT}�w� -��@��QAm)E�EJZ���-P-F�QJ*��D����F�4(W�*��!jM7m
F�|�P-�W�\��ӽ��Ȕ���B�	��wE_��h�7����p@�FkS{?o�;�{�_|���1%�造�e!B�Xh�|���ɼq�3n�"�U�.�6m"�[\Xdwt��[${դH}rK'��
D�����Џ����G�3%�o����{8���D܁Fm������nI��a�aE���'�{�ݔhU)�(���V�4��c\�%TiV��j��ݗ�goa�������B���u��"nkS4צ�>�Ow�z���\cr�D�Q��f���0��J2gGn�R���&�T���4�n��ʫ"�,�70�j�F�gL�n��3�ƚ�t��fjq���r��,�ً���~�'��\ɒ.�CaPxL1�F�ue��X�d5�C$�����l����CT����p�6��ni^��_�"��D��\m���A fA�o���H?�z4݊'N���VcV����|lu�	�|Vj��d���HW"�xzO��|��TϮ��u�N8�c[@ƿ'���UT�8�Lvщ�i���u�>?;ho5��4��	F �_6оKKh���q����\h�GB#@ Ƅ�Щ�`!���F�b@��j4�J4$�I6�	�24�i6FT�(�ڪ�Q���2��j�jJ�ibTJRBJZ.JU�c+�lDP�M��5�+�(H����o�Y�ܮ嗺�m��mF������o��+v�ݐuG��y�y��ei�FV�Xv��|ƻ礼�������k�x�z��iZT�'�#��~g��/y��ؖ���C�e�$z�F�R�_w�����MS8:c�e�!T�U6C+4C불G���kh���=�VԌ$���'߿qr��Vg-���6J�v���rYkn��	X<6�,F�c��*9mG=����맻��
��3#z|��ngz̅XS�ʌK��A����2�e��E�F�
�e�{�K��?��r�f�"���������P��6k��tP� ^��m:�B��f�i�5��fLX��E�y�qƃ�pm��|}��~v��������WR���>�ٹ̟wx����??�r
QC"5 @b�"؋,}��vl_�����Vl��㍅���fy����z�}�^l�>���Z�����_{W��q��_�5�D���d�3���� �bHҲ���5���uܙzֹBJ�.� �����EƔR����({M�-0�|�%0\� ^��g�O>~�ƿ>���S��]�Vf��FW0����m*g�j2͒.�F˕��q5s\,IQ�ۖ*|\��[%�g�(?`p���5��&�Q{:�uk��,��i��C4#
� Ŭ��?Y�<��f&��%2�ω�r�;�}����Ǆ���X��Ođ�x����F>��������!� �ral�#��$q��=S[5F��^��SG`l ,�l�A�Al��^-S��h}
	�n"�Np�l%����~~�8�Y�sF������_���j����F��߻I-m`���b$�`ĚJ�4W6�δ9L�#e���m��|�F�{ڈW����5y����y�keΐ�q�z-�C#�w����kZ�7y���/u!�c��{��}댛�&/�=���E��G�-Rҷ*4<�}qAWR�ﳙ��ڐ��}��7a��6Z��Xh�WY�R��i��i�m�Y^SXUNy�+f����5!�Hه��YR˫-K��uu8R�T���\@)�ك�4�%[�9�V�Kpaw9�:�e���Y�6&�Wc�br$i����vh�Ge�ċ��F�2�F�sYv훅W8#9K":�LL�k�l5��k�H��3�����k�b��.�FD��9�0�����F���
au�q��T�B��[]A2x���:.�3�}���|XT����%J�D��y#�KCU^;�pk��T�X�<b/,ڣ�ᬪ�>��ls�3(0�顋ܫ���܄+*�ܓa�=;^����o(�Ҥ�`ӊ4M�����-	H5Pe�����3� �����l�D�R(�P[+D�6EF�Y,��8X_+�1�ڼ�"J0�r����2�$�!-OY���qn̶�,I�ǨOO}݇_���y��/�ћ���?�~�q�$�D���Ĺ|�*i�M*�d��{���(?����ǹ��bB�1ދ��{��ŀ)�_�B7QN�|�;T襡EV�d�Ջ�����u�A�C���]�n��s56u,G�5���4�Q� )5�@�����֚�9�mTJ�nHb��0�R�q��mJ�`[xR_ąz����� �vK<���7�?g��*������gܼ�*P�KĨ�Ƃ ��;�UY�Mїl�23�E���d�W_ߙ�h�/ߤ���)�×���o��m�̈���S>��A��!o�Q�"���T��������h�"(����2�c[<�q'�Q7��4,��8��̇']���&wI�"4��U��l��{.JN��c�{Ł	6b|f�$���V|��}�7��3÷uOu�.��gփˢ�u`�9�4<���H�X��_kUT��-�n��k�g*�1QR�QTrs_n��N��֦����$���g�ݭ��k<���sH"(/�J//qs|;����B��;���8�H�f�ezR3��aMLу]*�^�E�+m��s�շe@ƌ�Z���H�f�p�||�/��P��v3�s�?8�8V6�h�C�1�<9cE����xc����)�/�H����K��d��}u|���{���M���o�N�++���{��=�?��r#�6�QH��4�����o[H�G`�sv�^tY�{+J��F���[.ţ����>��5�y���w�P��B����Ng	!��gg,Jy��a�Xp{����l��z[�fd��Bt����
l�dppv;x�lDzNR1wRh�`�b�����f,;�}����Ł�0w��}�t��K�?A{���t�FV����Ws�L��T����o�۝����BoD9|v�*/��o�擳�-�wz�{3��iۭga��̢zf?g�ͼy�z�ܐi�7�oo�Qnhڢ+�=��e�b�M�Al����2���gȌ�[��Z�s���y��|�I�]	�V2��������,1�
����)��52��_�=��~�.�W��~tjU.)UEmᙆ ��!s+��2��kc���'�H�3�f��CB*�@�)0	\�5<7����-�#����;Xl�z�a
��y�qØ!fCL�r%'�Xp����*�il�S����y�
�q������D�U��˯{�<=�Rm�I"T����y`I�$וz�$�"L������o�r$���$���fD(S(E3�U�ի_�E��d�g�gy���Uh�
�R�"0ԈmSQ������P�c�%�hu�+iQ�F�	pSn��R��(HJ5k��F����5�D�&4����i�y_5�Ǘ=�ӍW��rm2�Ji�F��[n����Z�*���_zSI@��my������o������F�$0ߛ�1��E���$�&ܒ����mW�/�y	���V��Ivs��Y���UƌK���u/J�^��q����=e_a�'��B��kxii39f�*�Y}�]�]�&&��QS��ki�˿������g��o��F���9i�^��$��������:fV�z�=O��T-/Oi��{H�N��	�(���}"sr�x��ٹ �d�(B��\�\*�@~Q� �槦$���2,ௌ�R�<�!ޘx)���'��)��ʵ`�����G����"�Hh���3�'T6��|R渙���A ������9�z�w����ZF���QW�:����~=��k��i�ۜ�6��+�o�̛ywz��U�HT�ҩ�&X+�	�o&qI � �Y�}��%�n��LY	|��K쑈ӗgg'ؖ]�K�� �$�x�,c�p�-pj�2T�i�1[ói��ɉ~%�7�yﾼ^�D�3�\���Ge˅O'�J,4VD���Zq�؞��U�;����?#䌥��.D�H�l��R3��V�j��CiҌ���*[�h g��WN�cF�&�cҊb�j ��R�zM��T���\��d�g���H0�׭��O�i�D�ʭ�؃=�7�D��0x*�V�B�1�/ÅO�)�6����	��C3��zy��y$p �PB��1�\l��B�����#���'����&4	ʭ�S�e�$��C�u���ii�6�a���戻`����!6t�7z*��P�E�=0w����֚�-8�M!YN�s\��o�����MA�P��11, Ҩ1>X�ik�ܒ��N��#���G]ȣ������*��r�Jd�B��ĴҜ����<�Q8R��f��g��C���Hĳ��&�ZF��S��b&��|}���|��t�<je�Z��+��Yr�d�t��"�ʕ)b�����W-a���K[���8 N��G����ؑo{��Gb�Z��L�Nyr��d(��C���˖�]�nI����^AA@P>7��7u>}ss�������
^��u���
ą���L�Ы,U޺��O�=�C����_��y�9��TP8^��2�Z��aX��%��N1Y��x��]�5���#��Xɥ��5Ϥ��=��Mg>�ޫ�R��7*�i���{�͌�n�}I��wE�򊭽�%V����^���z.�=�q퓞ʯ���f�]n��0w�	2W#�����Ͽes�Q�V�l�p��~��Yݮ*���F�ǾQ�귯K��c�_���:�3<<�c3�Pd�k��>8��f�E��
��_Ju�v��;�rĔ��e�_�7u��
��䚏km �|V> Ɔ0(R���<�5QQ�4���nZ�N���R��WF
���疾�`岤�U���" >��m���Dkv}ڌ3lD6�Z��0���Ú�K@�T����(�YV�"Ҋ�дB��^������F葋��7A��8�d���Ef�AyHl��[4
鄭�`���M�Vi� �]�-����DjLP�Rme��)�#muH�)��utɬi\r�Jnsa+�
�˥M���PꅸFŊփIFbղ�l�͕i-HJ8n��KrZLD.�h�c����3@k���n��x���e��au�!�QYc�nyVg���Yp�4����蔔�wK�&o^�#c��]���ֵea`�]������|.'��5�
L�,��wuc��;�p��Ð�př;�㢁Q1���4���D{z0<J{���NB�=d �s�ږ��ذg�`�Ҧϋ����;oR˙����R��NJL��A�w�Mj緙��~cX ���UA�GJ��t8� �,��V���H���6����d�[_��i��4lr����q�lo��a0)˧A� ���U�*^G��<�L�A5(=�N�B�M�"��)����-��;�:��5&$ΌfgN]�8D�d�u�u�[�,I�(�Ji,��IS$@Z)��F�m����9���^Y�F�z>�f�.��i�sA�X�"7;d���C{�I���h]rkvv`�w'%ّ��Vf��*�D�Pi���+z�^�[�ȧ�〳f���Yg��7�!�uK9Y�\�؃����V���w^fAłˬs4-�(���b��V�,��������A)��Һ��0�D���6qi<6��?���d󗽩5g�=�!Ri?s�7���w����yw����ϿߔY�I��Tm�?:����-�B}�衻*��+"����M��3;Vw�7��P�_�Ӵ���Rdǰ�c�O�w��{w}&~�x��Y��7�s��5ƌdb�������O���g�6�H��������jr��Np��)��Y���Haȉ�6�[�����Yg��>�z�}޿{�F+)0�	X8�p��!����$��G�7��� >���mLa3�$ I����+�-�L#$��M�^�o���ͭ�i42�m��zx��g�(�����MLoYsr�i2�ݲ/�A��	��~��	��tX�b�
m��:%��={�swL�+�(���SYa�A�&(���6�^2
�pr��S�3�ڣف����\v�����&jv�F�W]3�̴�k��΢kF]�sѹT���崃6���̷xCƏ��r�k��9`�K ��3��A�B!7=ٶ���+_Ā���:v�d��V=X@zcA�d���%���>����7q&��*=�ο����_�����^�87�e�d�,���|ޒݵ>�����t��2�;6\����f��)sb`�݊E�t�^����4��C	wQ�L��n�z����4yi��
ͶAꍻk��+D-��q�Z�>���:�sSvϬ�ZF���QP�B(�����L>��U�i>���	#�L� �:��t&��-��ҽ_��]���~�=���Sڹv�Vm���g>����~k_��nDhD�z��6�x���3��6��� ���gQ[KZdUc}2��az�%_	ʁ�4e������H\�F��8�=Cc턀@�yڹA�oC�����QI�B���\wK��1�� �E繻��>K<�>~=��?op��5W]���:��6BY-�)����L�v�a�l
�r�Mw���4S�hm6X����f���Yc�����
(��O��w����c̐�l�x�u{y� ��$	��+_�3�t/���ĊO�����[��6��u-Q�0����aEg7���g��@�
�����a${1�a!I�x<U�lSM���G��'�r��S���L�̎g�j|� %^�><��b��1��$�T�#B�h��Xt_�~�w��Α𢴋@~Դ�����B��(��Z�ۢ6ugy39vN̊wvv(��㶝��=q�B�e��A-"�oMP6�Xw>�X�W?PO09ax<3����$їuR�m�֍^
�Z�+a�T{r���ղ0_��p*��c�ٽ�p���f��皮�q�^h��U��(}Mbe�0%l�P�5�;��ܳ]3�b(;x�d'uN*Σ��+�QP��j�1ݚ��M�jdDs"[��.v���ZE����,��ݙ�&G�W��]T��v�ڑ������Ó�����}�>R��Lb�QW{���}>kz��������~-�ǹ/��5�65���;�w�Q�
5}�+��E����8����r�3�L�,[X-���n�uH�`�H��D@�tSƋ�ǃy̐�����5D������k�G����X�v`�"ʫ��S�+�Ӥ6����O,!�������Ɔ�heDػ��#�6�{�-%fAi�{$w�
���d�	T/��vvLć2H_hƍ����������b��$-��3O�X�`�7�b�E�;���J<�g��>�ɲk�Ɔ�1�+4�p�w��H��@��;�K��G�ZJ ڃ��v�����{zM
�Z��^nxTD�\l:�
)hfy��'7:t>�!�0��*]�/�5y3�L=��p�>:Qs�1��(�5�=5nk�Ve�ks��q�'��6Hҏ�Ti�hDH��m�� bqV��>y�����2DB h鳒��f�+Hl4����r�K����)�\�h�-m�m(�ʷ]ʵ��Yv�gCBb�˫.�ՉĢE����U���*�r-��M&1b$԰tvk�!t�ee��TRf�-��-Κ��f&�pe�ĥ�ܱe��V�%b.���:�IBc;JE��b�� MIYc�l�	]塩��0�ImH�f�|��y��[r��� �
J���\u���
�^q2��5�+����o��P�}�laa2��z��;ސ ���/��1�v��T�w�`�'���2����.�V�
c`7'q�51!�i���=R�0q��$��Ὺ��~m���9��B�� C �Xj������K�Ϊdy���6N,�}�*��#a�sũE���3
4~ھ��'A�O�_3��n\PӮ��\?Eic����lM�mў�ճ�Z$�����d�)�3GFqfe��$�p|�2#�D����fO�>}����S�>Ȗk�V�;-4���ˢ��<�%�x�)��l��:�䳖r����E�3 ���G�'d)��B�i$$<lc��k�eY!`xv��m�����xp�1��ϳ���TuZU�*�M�mt0U��B�vFW*p���\�Jfk�.&�?�X]�FO�h����`����W�pkS���AFZC�����O��4����w��|$}��f�7���^�D��~K���I�2(1(�/~~��Ƀ��*�8k�X�D�g�kB�4�D�P�O㧄'�؃����')'�ĥc��:ȋD��/�rR
��"1��{ֳ�-o�S�E�6���ײ�N`ZW���T����S�U�~�>w:x��ן����r
H�R��l����{4�A�i��i�����my �鿹�#ZB8���`�F�GF�|T�xH���h�|�G�ar6�?��D�I4�}��!g����&�y�<���~��w\�3O�t�ؐ�l� ���f�T����VK7���=��������ںa����w
d�,;&�\:p6��4@�-A��	�Ds"�FoZ�p㷋��YGG�ś��EsCܴ"mQ��S㿽���p>���̹�a5g%��J��6�[#�j�a�wCb�asfB,���|����XE��QJ�:F����^0��� B�i�|6�,@��\BE2�\�p������h��;vIUr�X��IJ���2��b�!�8n�p�@�lJ��Ì@Xu��N��g��{uM:Z�O���T>�~TBV��GtUS���j���c3�S3�8,'��� �����/͹����ċ��[���.o�k�Z[x�ʼF�٣pA�����N㦩�v���wt�6�0EE��;ݽ��j��|�p~���ȣ��Q��KS�?��k�$M��B��������>#��$Ų�0$�CӋ8�y��p|{�6��$<���"϶_S�A/	z����]�p��;:,��Ǵ'�˃�r�Ac8�dV�=�b�.�b>����=tf�Q}�}%��80�,z����Ϗ�/��1�1�1��[Wb��5r�*]�`n�"�m�X�k�b4�<)f�(�S��4cc8d<���ЯH��S�R�ye^���O�5*����ٱ=�8
f2d-6�rB��G�]���c̴�U���M7q,�O��7�A���q]��K�=e���2��2�gIԼr:�>�5��Ti�4
+!BB��#�!��^x˙�hVB$��	Q��^%�����&�~��Z�T�Ý/3x�|�|��+ʮ�*�K�wBG��Pfs���^FJ��:r#�9Tk�3G���*��k]�8���.��5�:��n��r�"�QO�{�Z���p6ce��ʃ9�W)6��{iMH*���-TfJ�"z��ki<H*
�x��,C$A��M'���s%lOٻ�~ʻ��I
�Y�~�`���ߘ�8�{7道$�����9|��XtF�m&��?S�����Ip��>��<M�:��{�����R��=�Ñ�l�2�2º.��rʱ����Z��s0\cJ͛h�~t��瞨�K�`K1wL���qC1�ĳ������acy�ho5!x�MW�,��f��S!�9z�Yߜ���!�0��O�3{��2\��7��lO5����{��a��1	r᧭�IG����Ԝ/H>�XyH��ED�M�BPu�ThQK�#_z�M�r���Ed��r2�5�F>���z�#�'�A�ko�m�g	�����5{Wx�dd��L�n2��Z}r�N)]>��)�lq�wN�,�;3�r��E���w�oչ3����4�l�3!f���Fd�r���4?�����t؝�E��0�b�-�݊p\/;�%x�L"�;�B�d�R�Si6�3�D9ø��赾��U�zf�ʊ�S����hI�qo�i�kd!������;TǤ�q��D�*��>=^��ib��7t(�+�ym/˟���o��r�N�sL�{Vno�',���=���XǗ�eW��m	�];+��u��0�;���x-5e�2@���w�q�{���ӻ��5�xN�y齛w��(D���r�{)��ݫ]���3�_b�{��Ӟ\r��0s��Ǜ���L��ئ��r?gx�q�_�qz)m�ލ��*��	�/���ǥ�^\�A�����G%�� �ݝs�
��-��8Oy��J�M[��m$���s�`�.�ve�}�;�w}M,���4z�����ST���u�b4�ҩS��MŌȩ̶%N�N� �rh&�dN�������3D�O�26�K)�`�қH�S�{,�j3'��6{�P���͈��7&o�f�
'پΞ#���=�5�g�oW�O
,w���{�㾅�\�ڮH6�̲���*�[U9ªI�aQ2v��fa�p?;ԑ���fv-P�9�o{����u��n�=�xjʒۚ�i�5�#Jo�K��a�,���E�^���ڧmu�Q�Z�1�P����Y�t�wW���ȃ��r�^���|�5)st��$��{;/ǌҬ��{��p��﫜
���5ᩤ�Yw+�}�8�f+;N��]g��\���8=O��{�g�fϵ�Oi�CY��?���ҳ���{F�g&�g�r�5k��#w�y!�];;�F�8��K�G�3x5���6����ڧK�h��zG|�vB���}us��x|}�wml�l���d�ٰ�U��㘪��R/��䬝�o��Ap�`�=\^�!��G����!�S������.I�6�\��!>;����5O<���<x'�G��@�����7�l�K�Og�v��ǹ�܂�fW��4�������%��c�!�i0�l�m5������W(l��M���r7R޲����ѣ���:���v�7���hcd��Q��L�+fL(�-�5�Dh$$ƉCJ�����id\�tf�6�/�vB�FR�ML1*hQ%��\T-˵��4�oVT;Lcu�a�cF6�8�;]ā��!{e�JG�����&5�M
Fj�e�w&GB��ٮΕ ���4��"�j!2���K���,�\$�	���R�ˌ�V�aҵ��f8�w
0�L�Ƙ��6�ƌf�n�3�B+���Ғ��1W[ΫX[��v�#�CLW,%���%Le���L͈��]��h�,�ɚJ4�A�%-��f�)X�ѯ!V6��[�^��W1�+��66���m[�
�0%���ЊM
ത����0��<-rJQ"����ۖ#�u5�Gf�8��e۬<_-��T�+e��SX��:]X3&	��6�5��U���i����Hl1�5�CJ�33K��A��d�E���εq�ʃuѶ!��5-�X�*͜�	k����Iut��(�h^S�.-L��0,.���ңV�6�h`�R��Z1Ik�u��Ј`pA4s�i�0u:����W�Ur�i�8�ur��L-��5؈V,u�W�GP&����Жf�2��u�5nz��#7`4S��J�ŹL�k��:i�0�9�R1�w��� j�l5k0�q��K%N�E�*<��1��]�B�Z�n�l�0�a��c[4�k[C.D�`��H��KBU�eh�.�4֬Ƚ��p���r�eir��4:mx�6��jʒ�[2A�p�!l8ZrB�l����:���-�Vj�c�P�;:�k�K(Y�u�XYt%Y�B�Kkm�Yz� ���[����Y��+n�%��oY\��\A�k�K#�Ė$� �YM��s��Y���K�v�=!T+�oE-%�l8�ڰfX�f
�p�.�)��i�6c��Z.F��R�XM�-GF,�@�WQ �z�,���,�¦Va��F!>�̙ }T� Wv�,��Iq�	��a�i�b=Fin���1���f�(�Oq�wU��e�_
�G�I��
�*a~�Զ�HR���p5.8��!{^O��Ɖ�B����k�j���^_�G�Iye�$г9�(3H��� �	��{c�g�8�v�6H|��&��b꿈��>X��}T~(�����*�VU
H$�c�"?w���@�Y�t���X+��O�4�n�W�U=�#���Q����P�Lu��2�Fb�"��w?RFaj�	!�aIt+���*�Wc-咬q����F�����FPK�g_�5�fnQ�7B,dD��Ŗ�/�R'�r��aCm���<iQC"Sf]e�ȈWGE֕�Y���p��t�n�2�Q�c��iC��CM����-��p�K��0\]��(�M��"YkRm��m3��Q@�L0�4C�q�j�dԘ�%���6vb�P�ս�1̶��s��H�U/1���ne%Ú�3.GQ�e���3jبR�1,�k�ve�#6r��nLB��T�A�e�`��a�gU$r�Y�@�ӽ��Y��j�ًajٳ/o�!.�F�0n%�R�$xc�ԕ6n���*�7B���4\T]=�W�e��_�����H��a��Ҽ�h,��
���~L4�@����K�]�؆}�Ԫ%�3|I0RCj5#��R�Q���D�8�(���B��чC|~v�@N+8#^��Z�V�
�--*ֳz��š��t����\{Yv�H\KӸ�v��T���O��\Y`D�d�G�.F௎0�D�9����:夗�g�|�y�ԗ+����7Jm����ׄ�;ֶ�b�&�>W�7F������[]Я�<'��rlp���]�8# �����/���cl��]��xO��^<f�@L���NΈ�ed�<	�H"`W��a�<����<!Ʌɨ{ľ``�i���F����$���ȳ�#�\�2�2uZFmm&1������Z���&�A�J���vhw�}>��~}X}������@�H6�Α"=��!l��^:�_!?��dq� �8�DK#�'��\�fV�I�~>��~�O?~I�����;�|��(�Ս�q�n7Qx�����N����T[�(� �H{��E���P��m;e�	$�n����z;j�g�s��IyT@�
Y��"">u��7H�ͳ�����%�;�Ǧ��3�,���w�T�x�@�;����I[��4��-�5���p ����Y�v0f��|�TQ��7̭VZҍo��U~Lާ��3�uF���!}��{W�w�sƽZ}A���ѓ#X9z�'�uR�R�ܩ#��GZd��{Y3јw�-��V���K5��q��N����Ҵ�|�!�������C���#��V�?�~ݬ��SI��f[))#N��!4٘����R�lv���"ͪ��v	�f7�Ŝ����;�*<$��W��ռ��p��3�5��՛��f�q�؆0��}��>/������;�}YD&t����n[=o�c�}����|c<��43\��{³JB��jб����b����Z3^�`>���{�D@�x�s�5�QE��Th��@���r����$̙�&vv���"ϤEvh�P�M��5k%y�^�25Z�0�[V�o����C`������k�5��Qٙ���h�h�pV���3(��Q����ENBR4�Ϸ�^B�ZJih��愈�4()k"�$�F�6�M6�|�c^��&�w����N�rH;��$G��㪙���P��F��YP���łM�>��is3�,��(X.�~)��GJ���x����_~���,��>�*�AM�i�{�:������~}�G��4;�6�NfW.�Є��x����ˠ�f]j�G�"�������f� B��e��S�vő1��`S;;;�E�D8s�c�0�uLLM�x@٫�l.���9�i\8V�J�}�:E\�[JFJ�3r�={�����!bT�C9
2�'Z�C
\�Ra=��� �5{�BC�W���y�(�&n~����f�ZQk�|'���O�����땫�4������>6���>���A�s���շG~*��/<�Y��j�<���=��(��]�N.{���������Љ˗�O/�����d�	!�sV�h�D{���$���l��>�y�5|����h���Y�����1Le�a�]Z��[��vn��f��!�{�>.�8�u��9��&BP�NE�t�p��(넫r9���uvo��2�߯������������y�f�}��l�i���<�U܈������䔚%ܥ�Ílj�ZTj�A�1���H\��ͼ65O�!78��^��k��>w��ORJ��|�d�u7��^ֲ4� ���a+�X���hW�^`a��:N��x;`���>�Q���3{�}��b}�A[��U�и�cmq�u��3ڵ��I�Qc��,����O�)��(��fhC\"��uo�c�����ѵ���UR�����O0�������r(j8��6Gp}�ި-��XY�ʒԔ]�����;�+��&|a�:���cM��!6�!�K%\,��k�f�3e�.����\:�0�͗plkR�l�FX���;\S5�v.�1pȥ�`�ѺéEK3/S��Ε�w����3֊@�������/|sP񱶆�i���eK���b��C}�f�Lk���e��~���;X��	 _:P�#�g�?��Ki�A��
"�n�K��`�ڑQ͵��Aׯ�ۖ��v���m��gϷ�/��2�AM)7�z��޿�A�4T�0٩�{���jcR1�k		�<�χ�"2^G��q��.D����Gu&O9UQׄ��}�h׺�Z�!�wH�2 mj��tTy��6��iU[(}��5���f��5��:],]u�e�se�Ф0Š��v��P�X��ƅ+V��h�����]p��pPr� +��ó	���&��^Ÿ,��gViXB�M��nIf��c�mL��eu�t�d)GD4�ʲ��dG������f4"5hB�a��0Q�[]�XE�eh�9���#oH���W6ܖ�rR�Ll�:].���O��Ѷ^���0�F��)j�JR��Q�+v��f��hU��i�4r)�5v��O<q��\���H���&��[w�pd��gf0(�|Ck��6Y�P4X%�u*QjBA{�~:��hg'���K���Ċ�v��fww/>ǩ��'5��W�w�o3i�ZU"(�K�Pb(����6!U�IG���Û�T��?���z�2��4���7@=@���;���������0�5�"2Q�h��o1�B�ʲ/��K/Z�n�>m e���ũ�&��F���J�0�8\��Dwf��]�^��U�����=|U[-:,��ĥD�qJ8�%�N�FЧ�F�)�5N* �=�s�+$��ܢ�+I;�1Aٙ���P�V��:��s}�z����L�5�7X�����Cq��w��=�����~�vEl1H�\�&�,�Ҝ���ј�VdҢkko�T��[��Ӌ�%�aJJ�p�K'�T�s�-�Zm�k�&TaІe��ǀe�����?��Ę��~�о2\��-:t�D셄n����UL�)F��Q�og�[�O_O���[*�MY���z_�k�=����px�Z��EԆJ�(�#T�C�"R���дf����vTE�I�2F�|�bЁ��-W�A� �V��9r�ƀ)�����{fu��)���:�#-KH�F
`('�ʅ���d0�cxOo����k^�s�L�C@tn
���D��� 詣J7�O���w$���t8�Q'dٻ��݀� VtqL"h(�[�2��7F�� �(�-c����g��1G*+�9#�<�u�]J��c��]Ğd������n�n�Yb;؀��^�G�JMa���j�5�Vw;�~�x>�`�5��?^��j������T,�κQkP�:;AҢ���8��XKF����Aﾩ��|�R%��_a������@����!�F� �\u�!����i�)ˀ<H`Uy����Hİ���Ɵ��4q�Q!	R��a0e(gĒ# q�]t��ܪ�p��EETV@�r��|rs��g����9`�>pZ��[ݺ�ܓg=ٰF�kMa���=�v���.U�*�Hk�Vώ��Ͼ������(�g���8C�6�<����ً��h�i�T��4���h4M4��7�)��1�Su�zd�S7ͣ�@6lM��M�`��#�)�o,��a�Oezτ1�罻~o1�,�3-�n��w���[`6&�_=ϰ-������.��_ny%���P���뼣Mm�/KR.l@2U���Ö���;v+2�8e��_�v���#���x|T=!���ԭ��g�.$����b�š��f��]��ѯE��0a���X�3<ԯ�;�'`]˻;�t�ٕn���Ivv�m��J���Vh�*��a.E�_�;�_<%XQõO>��i�	���}<���ZgsĞ��YȏfA�>yύo�~Λ�B^��Y����y������u	y��:j��	WW*��1!�kg��E5��g�J;�惀��`��H_T�����/�Fu�O�>�ɿ��8�>ϙ}e��S����ULd)ev�N���?���%�����\Ј��oa۝'bl�'l��k/vJ6(�>Z�j�8��^"�Y}�s�\��Y9_��}���؜�O	^t��%��Q>0���˯ôSVc5�3y��[�؛獖�c0Z�C�4X5[�оw����PAD}���]*���=�O���1�Ir4�U�^�ss��8��^��~��*  -�8�i��A�g������>a���6cLp����_`_"0?Gh�6�W��#�Fi�(����1*Usl�j�5L}��U�����k7����ҟ}BU\����nƌ��d��a���5�`h���P ͂hca���_�>y2�e$�vD�F��TBڧ�-Ф:x���}���TiY0;^slX�zI I�3��m39u;��?l�J�X�w���u��b��L�Y��D��=\�ޛ@W�ZD�uv��ހ��2�p�}�h1O��SX�>-߿�����(/�������2D[�6c�y�N��|TA�5X�.�Y��(I�2u�.�ސ�,��q.��a��G���ʞ�c��`��i����`B"�i�>�����#k���=�����_쉌l!�F7O�^F���@�ű�p.F�F�<��v�h%�OIF��̖ԐH	I�C��@�;�3ߢe�|��i�p��+,�N{w�١�+Bm��|���DN�/W���w�"��p���e�Xv`˨�&C?���TM�Y�)�lm�J��E��=�mZ���o��}ZihJhG���D��#=�eE 1�0mW�{�H� F���a�v	�l�n�L��[B���:�,�0�k�@n�0e�8�SJ�(�ʺT���l��Z]�x��15�Юб�˦��J�2��X�vԘ*�X�B8v`Gb������87dA�Rl��-���j�k�����
뎹Ź�v�,��XG�̼�nּ�H�n�f�4K,���\M�:��KJ�Ρf������Kl�U ��6�UJ P�oI�!gu��K�z"���<r��U�V�a��B�,�6�$6�넨���I��dSYQIEv{�ߡ������y����aR{����տ��,׫��m1�%�E("l9��ESF�Z�1F�^��F�""�C9��r���vNY���p���z��"���#�m�����ۉ`�J�n��Ꞝ."6�ÑD�V�:%��86T���|g+�L������Ѧ�%{�k7�@{f":�1�����"C�͠��9ݱ��(��{g$��
�9.�&)8t�1}�.S��}�(i�nO����G�W�I+mZ��]0��=>���c��L(�QsmU�E���<�`�����jz���q��N=5��i���_l��83���#�7!��-�~>��y�P��� ��oO��������fi�p����#��M��ͬ��{ Aa��l�4J�
^:�BP�G�x[m�H`�.��P��R��r��֩fq��ml�3�� JBD�����:a̿{:��R��4B%-�R��:E�	�+��O�8��>Lk���A��]�-��l��A��Ԑ���U<�'}截}��a"��xh�#��ۏ/듷��]�������۷�|7&c{����ZB�2 ��#I6�Chm	���h#��T5�M��[g������1�0) ��Da=�q��XR�O�5��M$�w�J-��b3N��zOhB
�	s��� ���6�I�Q���E��N��N��U(��6#��>^cq���qc7ֽ�WX|*�ք`+�@ ��p��z�T!d�8�R,��#OP�00� �1�e�@�za+�>cDm(:�;�fvgN�U�i}�s&��}����a���Q<��:h���>�y����Բ��au�t��'����'���=�W�:_]3��X܃u ;��K�4Y�Z�00����[������P0�L2$	(�v�?$Ȁ�v�¶Z���A<b,*y�x�!�h[l�����UD��6�ZlQ�ƐcO����sCy�-�ѤE��]!�ȅE���un�����6�-��W�OfEi�4�����H���[�%&��Q�ٜ^�"��)>I ����Mu�:���`�x����߿a����3���?>�*lu�7!	r�h���;�a���m�k�X��v����2o�'.�a��g��&��ʹ�ͳ��
;��{����^�Q�l��F,���rr�M�t1����ƌ�&ɾ;���2.G�5�"�gnp;A�Æ_��gwy_������$ѹk=��NDvd��\�}��wt�_��lY���ʷ�ȐD����sS�}}߿R���t��{b^�<=b�6$��.�^I�� |���xf��U�)8�G�f�-�����ڐ��.n�E�7�	�3�������i����|9�˒��Ov����q�f��L�Bz�7}�X�X'V������ؼ}�;eG�yzH�l����{��oe����K�m�g��;��va���_��yy+��r��6xs�k�f��k����xO��]�S��a�{#�2������n�pȱ듹�8O��뙻�\)�S7��C��L�j�WR&$R�,�25�ʶ�ؘ���^�
�E�-�">�vt��}Ỽ'ۯ�,�h􆮠�b��&@^��(��H!!YY�]�shd`�Fbx=���O�@Z�2S��u6��i'u3mxi�e'�(�{�F%>ד(Q*�n�w�$`�'`BdE|�#�<�0q���{���Xc$[�啜ɛ�l�5��	��	��+A ���+1���1.��p�&�� ۙș|q�5�:~��-�|�D�3Uv�p�;�T�ٚ����ة?�*ְ�H��?��hqo1�OǢ�?N�ٍ^����`s�{ۄc�]P�6Jğ�&Ao<W|���N��۠�kj��V��Pl���������	(�s۾��@��,|[2���st0�G6�_�/�t����%/�&B��K��4D���D�A�AT]�{��"4�!9^$6��u~�Qf��U���2�A�鞣��gb�o�6��\���4sZI�u�`��OCU���KA��]�o��y�auش��.-;����Ƈq`��P�jKdr�heB�,�L5��!R}g
��J3k���'����+؛�2�!��17��BM<�2��X�\�w�`��ҋ�M`��
f4qq���ˌ`}q���gΦ���]�r]���/���a��?c�{��u`�1������ʭ=(� mH4��6[@�Ă4� ��r2��G�����f��t�������4ES��m�8��"��
��wzp>�3�ܳǦ���9+�>dχL�����q@�^vZO�x���FӏC���Z�3��ߘ�qU��&�M<���9�KIр^�`D,T5�-�k�v[q�GI12�|��\�B5nN�Us�|�=P�}dnO ��ŋ�.�!���C>�j3�Z7*h�Ʊ2��^t.���4�����&c�ΆfH�ɒ�%��!����q��qX������^K�Lb��Th~��߿~���o��M("�!p���>M������{l�>n�����j�5jF�fx�-�bݨ�iY�t���_�z qQ�U�/��6Q|9��cw���rސga&Hs5������n�S�䫸<e���)cNɡ�2}���Zl2���]���@�}��� hv�G�g����o�;�����=�)ƖQj�O�C ~����e�
b0ё�#�7�j�0�r����	, �G��>�NT�f��%�pp���l�_����E��B�Z'�*pF�J*��+N��"�M�|��>�U@TZhi�x��:�R5��������TTAJGp$�*ܭ5�ўC���~!��a�r!������{����5T�>&�����:5�1�0FZs�3y8�c�W��G���UɀN�g=O��焰`1������l�=��	�s�\�������R�SS,.��՚�"�b���&m�d�3L��%�%�K~9��}_9.�Z�»����h���?n~�~�;Ki��_	����v"q�d�w~�Ӵ�q����<T󤓧vL̝;��#�i��4h��-<�iU�v���>'�C�O���VD
LB�f�ð ���V݉�~`t+���p���ňw�xH�I/#�>�ZCRl'���>��?X�?�n�}��W�bu�>�"*��| 	"��3Ǌn!rH�b�2|o:��! X�C��5q��s���
�6�s�s4U^��ʂ=g0gt��=ߛ����S3s��9vgI�4:�gq��匚�9� ��$�h��͊ ꄗ@��Ctf��D
>�ZB�y���&�,D(���ڂ��x;��#�c������h��D�9��n'LӨ��
����zS��JiA�����YqI�>;�N	R(�wb���c]�r��O(SxF,����j5��T�)(ц���e�X�� ��X���!����jg=��v��1�a�^аt7X	f��r�f�@v���ݰ�,S.��N�B�+��YW(�\5-�`�wa�fC%�2�e�ƞy�g[���\�ƍK	xh�5X�%��75��^pؽU�KTњ��q���#�]�ڱ�izz�޲��%(��J�hUQAiDV�$�D+n(��j̻��\b��ZfE�!p�6cef�h]�����Qt�e���UEGbf8Dm6
�1�3��{�|/'�jҐ��)YI�(�
�өz<Yx����\q�`�#WSS3�L��d�3@�_�ʐ����a�k���.�W/e�舌��D���8Bu_�Jf锣�mq
��hh��zgyKkQ�jE���R:`/F~P}�W����i�W qr5����Ɵ~TD��9Ǔ�u�4~�����뎇�~?��(\$�fZ���!��Nvc+�i�g��B�!2��z����s��oʑ4w���g.I��%��(��WF�)0��\�ߑ'��m�ڵF��|߸��Qf�ڳ&�q��esݯo~vfڃ�s�]zD��E����CM=}��Ռ�YAj�\<�t��yj�e��ں�� l�;u���h�H�&T�ff'���*(�~�Lu5��'#9ʑS������i�{z�9����8ZޖT��gh��A�*�3R?�!���3f�=Ϟ\u)��C��5�f����e7@ˈ�K!�V^e����,��F6F",��yqp��w�w��������~�qi�Dk�&��f^�ﶱ��;��m$�Q���j��~8!-ԓL(��)�鷆��S�
Ґ�<O'ӵ��	�_�����I�ˮN��Q:j`��t$}�3��tj}���;�����O[���N�����{[��A�+����&vvI�G�J�O������ S�҄�����3]��bk5��:;�\iD!;X۝��CA���LE�cu8.�vt��gL�U
�ԇR9'����%��8㚰���@ph��Z���։��vq?~{��'�}a���QYi�y�͑!C�P�T�U�S��\��4��`%]v�*m�`��:0�fwW$�y�˝6m�x�.����^\W6��#�-���M�0�a�_R�؍v�xz�f��C�N.xw�w��)��}�gfd���6I#�}N��)�������u�MO[y�mй��R���5헸\��pB}��"�F�(�9��ݙ��tG�:��D�RӺ��h��5���i�p\>>6>���}k���{�Q�uq!=�x�wv4:��u�Z��mm��13����[O� �A"5^J4�҆\;�M�5N�V��Q�P�%�DE
Z�Q635&Ì���D�/r����c
jon̖'���,*P����N�GM1m�>��`>C�C;�\ǆ���3Ex0�V�[l?r�:�0e�"��	F��{��׋	�e��#����6k3��}��	��ZO-v��F�
=�H^z�P������uܝ�	��R	W�`w{�_kQn�(6ҔG��=�S]T��ZE�8�,��+��s��ۄ�3lg<�%���u�̴��M�=��1���Z;қF�p�k4�y�@�6���7d��V��P>�Q������A�z�K=i~����?~������*ig�.��h��|(���UD�l!��mJ,0/(H�W�t���$qq�7��!��1��8�4`ЍP�lj��/��)"�����/U&joY��l������՗��g�7��2��k#s$F�n��HA!�!�R��
~-�����@���Q�� O}�'��`���uM�˾�s��������5����-�huiFPc�rL,�yZ�Jy8�rs;�� �7�&ѶU�4�j�V��ɆW�%q�`�����xda��1�JL`�����a{��CN�$Ξ$�m�u�!\=�x#���Z�Ax`:��0�籖МI��=z�gg6�a���6��oB�]L�¶Xډ�Iy+F8�&�k-��2tId�f�β�Pɀê��`� �l(��eY�"�N�%�hh�κ�ǁ�E�Đ�.\�p��>�o�ѕ������}�g|~�|��3�}��װؤ7��F����D�l!��Ћ:�#���1ג���Vf�nwz�{����=@gv���]��i@ʮи8��ULa{��gǹ�{���W��I�_�g}kD���3i�������x�v9��}ň�(
|H�0m��AH!��b�����Ʈ����I0�^��������_~�f2����}|"��O��+�dzce�|�96ؕ��s���u����|W7lHX
<-��Ã1:@灈�Lh���{�.r���ͫ��=3�H�H��DE�]��t[���l�<I�
��q
��t˫J�����ݧ����Z�S4&�R���\B^�LͰ�A�%�WZM�K���K�G
��:��\e��"����WKՎٕe)��P�q��R��՚��t�BƎ)�� �Cf�-�s�tv[a]e��R���h��	������"v�0���(fX٦�����"�f�MXJÅ�\�Y�$c5�s,Уj�+6��*k�D��)\`�3�2L>�4m)J�T"u0�i�ѭtU�,Y]�h��mں�6���+j�宬�f�fJD�`�����V�K�!�n���I����h�ұ!���)��Q ���2� �H6�][{���<;��,������9 ��#�x�����X!��q�=h���L<ʡ>x�d�:�a�������;P৶v208��/�@S	�`�)��K�)lH���q��}%�4�F��z�+3�U�IWQ�f-4٫��A�]�_[�A�H�Z��MxL�L1Eoj~��L1;�j��i����GFQ&�0&���Xm�k�O{�iă��d=< �d��l���+!�-�<T���t�2��E־���w=��ff�{�3������Bllc@£��z=��xv�@E[K�o_Oڽ�p�x�]���]�"˶��6A����9�t�1��\�`�ۉ{kY[��
���(�P�dv���u6���AZ}�fݜ/��u�L�+�@������G9eM��2��Ba���w��j�!1�F� Ⱦ�8"��x<�4�[\�l�!�R�/8!34�Ƕ��V�mlX�z�a����,���[�������>�v�*)Ju��]�Z�aaCL��g!A����-q0��#5L�����ka��H���n���T��;��EӔLy�@��9p�$����CK��z�m�H��_Ct:�n�b8=�E��O,\oMLa�����W�x��up���}~�v|����d�q���P��v�!� ʰF2|��y�2
��LGe0���C\i*|5s����-%����+]K��~�p�؏7����R�T�4�� ��2���85n�vQ��=5ȷ�L�/4P�Iף�,��9E��]��sD��ٴ#��LF"R������*݋[\֘5T�ZSk=��x~��%F�	�D9���[O*��9 �蘩�b޳Y�i���)�n���*��>p����w���^#�n�g���ڏ��E����.��-Jj�5�x����2͵���m�w	a}�i��-}��}fl~L��������R�wc�.��R�י�yJ5�ϧ��<Q5�Rú��2Mƹc���6&���P&Y�j��L=��8�R�4Tjl���o;s����Q�)�H���M"/iDDSnf�b}��\�S���.��tut+Q*$H�I���6{��a� �b��ʷm��떷[e��K�	0ѽv����ƐH�{�S �I� �S]n�P,�#c��۴�>��%w9��V�З�������!��$d( q����W���_�sȦ$�I�O�1{�w��o�((J��(�����?3[�_[f�3�#��_�c
����S~�!������_"M���5��[-��c)���iu�\�2� �n1Wk�eWl�;�<��)��2���`��qq����G	�	�bH4Z!Bꈛ+�ֵB�#Dm�lt��A(�i�I�9r�Y��'b���V��&gOQ�3t�Yy��ޞ̭v��o�eKf�e����][o	��E^�2t�~@��2AF5�8r�9p�K8)Ή[�\ϐ�3*`�9Kt��N��t� �/����gK(��x�3b�F���켹i!�?;��=]��NެG����r @}jy�4���z���
��i��⸶�*��A���n�X!�,eXaHdU5��f�7j,n�K����K�]����.�GhFo^�w���{��}��@�R�*������y�������M*�Sd���p��~!�猧����'vO��1���?�$�Ŷ�̮t��XQ�W�s	q��`lҽ}�����޼���v	�436�=u6닥P	^AJKiMYe�	]�j�!H�}��a_ܱ��\ke�z�Mz+*�9�ck�["�^�hN	J�[��u�N$6�R9�F<��������?��ؤԛ$o��- T��@��d�w�&ZRq%�s�UϤ��j˪�~ʫ�f�����\�mp�B,�$�PwF}!��w�Ht�6�iΪ.�xV�	=)�*8��mD��z���h���#4?�s����;���;�ۦO~�����1<!sH��,f�����$�lh�ط^�xu��l�eҍ4�4�(����l���"���軺.��%I���8t����Mj12��z/ �'N32le��z�(=�NkӽY�jO48����D�-x��$�{�	�V�m���;��D�7���n�Ǖ�=�v_��^�g5��}�z}z��vk��%�|���%G��Fl=^�w�ݏ����ޟm%���a;�}�8��}�_{�����OGK�eoM�6�!sk��z�c	 #��F��Pf��}佾�CSsQIJ�"�vu�
r�y2����0��A�f@��Qs>�#���<�p���|�y�Y_;�����M%�E�������ʬ�L@�x-kH�b�r��,({����[���Y3NzV��ŏ�Tԭ`+�]9Uw�6p���-WXS�3چ<�rն<T[�f�{Q���-�'���Z��&u�;�q���{��9����&��[Rq�eb������2or�a]��+��R����ӓ���To��`��`��YE̝�J���<���Z���n<��i�|��Zi��qc���G�d�q$���쁜,<ʥ��AD�X��(3�J�d�T!��m�he��+	o��(s޷��D���a!�u1S��
a�J����1\��4��l�Y8�sI��:�qղ���a�LdHDu<�Cs(A��V�T��7�2N�Z5�Z Q@��bg!���D������1s��͆(��v�1�wg�kJ�5X1��Gb��
��~��	(��rJ1/eh%�d,j�cVx4Oԓw��Yebx��C�]��12��KK�p��*r��rq,9,�eX3�e�T�dQf�o:��e�`k�M	�	"�)�V"�Ã����w&KZ�2�0��f�������)^\���2���,&��,fr&	5��`M��،l�#� ]q5���і�1{4�d%�^{@a�xb5v-!G:hu�Kr$ֺU�E8���E�@�"B(7mvf���ch2ٱ�A�.u^[eČ��%�e�c@p�-�����%�lA(eq�3dŻ�@2�]+�3�C]378@�#ְ��^\�QΚ!�F1�6���`ԅ�j.IE.�lS&�*q��n��Ĳ�r��i���\m�KH��h���ɩ5�K����P��S����ft۫JR�Pb��F�WZ-�R�K3Y��Ն���F��ۣ��m��K�i˳5ԍ�]u�5� ��B�B�	l�ʻ'9,tl\��]��&�s*�#��sL�����X�u�+�+�]V�5��%Gbؓ l��v���B�X[����4�Վ��@+S=X�a1F���K�eF5!JY4;M5�r`�q�[�Ms3�;Z�;8�W��Y���T71�iE5�62Cڑ]L�.�˨Qf��Q�����F�^�$�$Kr��+5��i\%����cK��]��&�� ZK��d��j��9��9�ZͩP�ô:ą��]i5�ģ����p.�����%��ͳ-.�vm��L��� d�e��QhEGK��l�&咵CT�:��qL�`z˚���X�Zuк�3rCm�9���F:,���`Z�\�e��Bbe��\i���a����ѳ3
��3r���)�����B7Z�Bڡ��5f&#�)��\qv۩)n��4��
�jR8���c$�.�6,R�F��%m���[x*P̦^(&7Z�m��1���9��`�R
7\��&lL�T8�#�
3�&Ŧ�4Jh�$�c+([�vH��f����),�r�́�ѵu�42�F�[
1��,5H�R��3X��8�	�B�"VUi�pIa-��o�P%�������������~�tD�b��l��<QYgz�C	�ϫNm�Hnrrj�0f!��r���>�8������ؿZN��V�Jv@L�:d��T
�&�&�TCx�i��Gopv��0�\%&�8�/*���Pe	R�!*�X�n�����y2�-�r�|�Л��|\�"0�Ӊ��#��t�o�gS=���B�)�Sknj
����XX?�?x.�N�f�o���J=! �`�	�:�?��g��,A����'�������|D�Be�cn�]�U�ԠB�<�&�-s����f��-���\��,�̶\�\.���qGPzX:R=a���Vc,���8a�{3y��m�c6b	��J㛩��$ɡ�Qڷ��![��Z ]4�X
(] ,2�h[��â�@�*�)�K	U�UW@�3ufa-���&Y�l��%F��ael�B�.#K��l�ǽ�t,��\IoץWe���GYc�p�c�Kfflv�5.�� P�I��kAٛ{�Yi	��^�0f-ݚ���߾�p}È>	��L{�w�D�����h��n<�f��UQ��[��3LĦp�ᘗv"�0<D����//	��l�Wd��$�46��2s�<���jQ��z�fg�M��=�dv���Y�����:��������Y?|��!<.��3ͺ�b�5�/�u	�;�d\D���Ⓚ�0:���ħ�Ƭ�X��m������O;�BL4�8=��H(�^G�Ky�����-�2��b�"��*��r�m��@)��Y�%��ǫ9�z��R8����H��Cct_���}D��[	�Pۗ�dc#���s��l�V�� Y��D���Ni��9t ��/gjȸ��k*Ĳ�lÁ)[U�L-�k
��r��y�xRl�])iq����oK�Z�p�����9�^1�$B:T�/!{���u����ք�3���r�$���xb�
!��E�����fMp�����'"C�*v��i���6��~�w����ݳ8_	B(Ƿ�"-:��ZZt�2Q����jP�H��sզ�Э-tAB�Br�ą�X&�6$Ow��5��y�8�{��Hx��aX��;�,&:��N���%)����r���'���f}.�kA+�C1��ߙb��Md��"�A ��o�C�<�����,�^nyAk��ӥR]�C��Ӕn���;2B��n}�=)"t5�⧉�A��ؗ��$�Z����}�C���;J�\<��h^�j:����FC,F���!�Y��L A���8#��6�jt��H�cT2:ĳ����3a�a��3��h��Z�ra��-v��mb�����=m���[\�KV͋�E��t#'����7�E�mb�:/CV�������}��H9{�%كQX�Ό��L�튛ݮ��݋���	���p�I�J~'�r}W3r������g��f�$h/(-��M��[�R��舠�t��E�,>�-��JI�8pY���� �n5�[Z�����9��~�_���n'A7�d��RF`����Gן��V�)Du"*(+�Q�i2�{����Ц�!_*�DA��5���a����,~7G��/;s���C�������A�
E�K1h��l�,�q@�\�0]D4k����2�I������e��������)��h�+$�Zi�F�0E��{����������8CPB�L�����Oh=��t�E�m�WD1`��RF��:D����fQ� ����rs�����Z���i�Kv��F�[�d�J�c��P�V��2:��+��V�3�?��
�mҸ�k�0��<�����(�����"�#z����:_��G!�2�!�2�<���~�R `��1��\�%����7C`k{�T�,�Z���rcw�2�������P"�q�!��CDv9��x�Lo*�W)�z��r����Q�W�A:���s'h��W�4s��fp�PF��7�
���`'��~TU�5oW���Ά�"4��ONW���`��2�1��#�B�EE���Ν�X�E��1��į��39��c������ktY��e���F�]�vI5A�yJ)j��� Z9��w�����]˳�&.�K:w�����'��v`��X����	�4{���lAw�$��BY:5��flI��l/E��&x��*L�qu���P�]G֕�cL[j n��uakvp���*����i��v� ��1�U�.)�:��a��>�1oo誒�˳�Gx ��2I|��.z�Yr�:�	����
8���q�>��т<���Wp��i�z��E`8%��BR���AE3�|�t2�m�T����#22�;%�* �O4j��4�:+�0�����g�������v�\Cϼ�j;b��+zb�u��@�ou�ف���%�N���5��6K��v�H�mӈ�9|����k~��n�����Y�y�;7�O m��ԗ��R�tJf�-�Y��f�w��osX{�
I��h{�	�ovt��9��.�>�[��� �L҉�������_� �����������u3�iyH�Z�9* �H��9r6�ɦ��,��Ik�>DHnX�h��L����My6��MA��ʡ�@�SmX��D
������s��+s�b�fbŎ�R̴���eф�m�).l�IH�vKi4�ƀR��ݣC[u�fiH�ڀ&MiB꺴��\�2fblP�B&�&vB�qu{�#����b� ��nԴıظ���q4�q������ ��n�u�2�9��eo7d�B5!J{�ސ$�)������w4w!�s\��.���6h�Z�9�dP�Y��kB�n-�@0Qn�%Y*�P��'/�0���Vɼ��rdrW�#�q�TH=�j�==^P�h�/Vo{侹�̲�,J�KAl���G>�*H�x.؅�lD�[�N��7'�rk[���c7����,�"f�i!�f�C��l$4D��EF�M�i���� �#9	�	c�c�"��A�12Z���Y��wweٮ�qϦr����������"��GП{�5���@����:�1��ԟw2嫞W��@t]��L�WM�H�lb�Jt�9`V-���GJ6��B��y��+����tܵ50�!�{�n��
k��������埶y����UhJ�3��v�J+����<H8p�M�.��$��K�q��~�����8�F�qx>���K[���P�ZF�v���^�߼������@\�&���(�1��h��N�ӗv����|5�[\=(|�-q���]��U;4�x5��<�!�HoZ���g^�m��"V�Hl���f�� ��A^Bd�nTEEF��풍5W�UM���4
~��K@���'ޮM�W��3�̈�J*,3�N��}_w֐�i����kP���|~���FU��q�r\[�1�zi����iu2ƾ;����]���Ϩ��(Hm�.(�aX�E�BZ⎐(�%���t�'rI`ƪK6��f���Ϩ�&�.�b)KJ�E=���Z��Ý��1�5�B�Ϣ_�����5�����kcO`���MM٘2L\!�3-��$^$@��!G�^Ťh��U�"z��t��)�	�O���"/_��H�[4u?���!��� �}`�8���&��\;32���q�Rc[H�bb��`q
\�u�PK�w$�:�!W���]=��)�4����2�k���wEv"��ėz���Ю�0�)8��b��h8�1���Q뿄p�b	�)4��f�����	>���� ����f�$�Cp�~!�{���״A����v����/��#lRgE�̂L�}����FGt��c"�^���,�y���$��:\�ʱuTm�I��GN3����{{���ؑR�y�y�O/��u���m�X0y��� r&��&��9�]�g
_5�tc���_���Fy1�H�
&`x�O�!�E|X���mZX0l����o5�H#ͽ�r�!B�C��\"�<F�6��P��Ȏ�yܬ��Y���s,�p���`�6�FO%�8�P8D�2����gzO��m�5~���(�Pvʸ�t�o�$y���;~�붾�ŋ�J&��+n�K�	�it�����^%r��k��9��جUڻ:E��!WO�<���=,\@A�m�Q�e|b��/���]
G~��Ko,�9�ݣ,��%�&��a��@(s73�p�����B�DI�@Ꞣ�]�&̋O�S�N�\�Q������*�0�vpsF�gpR"M	A���S�ΒgwE���Ѳθ:g�8�����g��iy��2�{�1@8�l��<���<Z5��V�@���5�߾�\U�Ra�W��N=s�y��Z{ihTTh�D+͚ۮҼh~S��ӗ^��G��3t�M;YvqZe.:ɬ�ʖ^i�j]�����sw&&�4\���6��W�V���|��UBV01�bGB�?I�3R̐Q�8�lu�@��C�(~	��^ߙ/�b'f,da�� ��z��Jg�pj|֥���|>U½~�'��-�g���z��}���F��@�Ub1~
,akP�]W[�3S�0"n2�6�V�ѣ��M����%x(�k�C8���|���s���������'G����=+��>ͦ�<�»����_�!@R�i������=������b��>���I�>S\�]�/�a{c
A���<K�>�n�(Tn�cW~�>�l<����}4z�9�'�sWEGe��*�����0maͮ�4O���O/Fܱ޴{�»���mA�i���{�S��3���V�E?|���2�,r]�M�-�>�;��{���Р�sI�������p��(��Scw���t���a6�bQq��Ugqf�gLR�s[%�2n�r�
ᕷ=�eu�L�W�gaz�	��},�O�1;z�����6�6Ǥ�(";�(�Z�G��W#���3��{,��]]�=�����O���f�<�&򸽪0ŀ�����Q�N�kޗJ*+Mu H��ñ
@���@^6�P�D,W�b�g2Y6XL����65�+8ѱ�ؗB�SB:��3vcF��l�1�ӑQ�X�r�M*5ʭ���X�@��M���W2��bjh��C*�du�k�f[�e�	�Lf�#���-��`��6^+��6
R��cEA5��n�!5p�\�%�3m�JPR�Q�7eSh�A�aԅ�*[KkMJ�6"�b�Z��	�'tǄ��ig���VͦLZ�.��V�%�:��c�5m��<ؓ3-��Z�
���Ě˚�q��������`�-Т����!�}uƳ��L/�ź���9K�l��k���f[ə�V���7g����Ot���_�g��7��f���I�B�{Pja�\C��X��>�g˱�
Yz���)#����3�Jt
XX
���0���bi�*=D0+t�1d��Q�$�RJ�������ٴ�á��Ci6�֩�s��O��ig�C����3c
e�쮆��1�A���]{O�'7ҹ���~��F�;��aH`P�^�z��s���<��C��@�q�p>cd_�Sgo����.�E�E\��:5���ޒ� l�O�&�f�O�H�"��!9�8����b::�R��pq����~��ߪ2�:8�n�1R�#v�8�ƺ�� �q)��M��3�s�Iv���&�G\S%U���Ã89�n�G�"���$��C��.#��b>O����~�h%�h����m��&�Y���gD;��dS&oT�I��}��*[��3nB�J�;\Z���0�T��wƦ��x8��x_�gvM�oo��{�ޛ�|�ZDu	��7�l-���N|siϦ�=�8vbu�#��a��ys4�X�і�7;��ӄ�$�#�xqeȳT��{��Aϕ���i�y��#�l��N��`G��Lgɛ�.��5�ӻ��ɲ�8+����H�p)���Y���.����uTp�m0/�<���!��D�l�K�qJ�B��b�q��{D	|�Ʒ*U�KB`Yc�͖�_�~�nI!�e�c������Ug��/�8�v�f��9�gR�YzA��d7��D{LY^�gu@�B�oiD�Sm���A���	�X.1(�[�j����%c6ʕ�6ј�sH6�K@��h]W��o0װ�������ĸ�L�Zf�oǵ,��z,d�O�6D��� RDoL�p��\���"��/X��Dt�$v[Y�P�g%�un��nIxׇl�t���o���ɧBt���n��K�\l��p����k$�f�5�e^���D�Yϯ�g������Ko�k�e�w�4����v���K�bCy�Pseխ�2N7�[���"�����		�
3:v@����`�8�ܤr�"�x��t.(5�E�J��K/��x�������C5�]\Ɖ��X�|��|��Y�5u�uy��Wh~Y3�:�Q)r�>��񇬋}؏����ݽ{��I��{}�~;�߲Q�K30���>�l��_[(����|�}��|"��Ӕ�S"K�|��ȶį"5����9�Y���1����@`F�1W�[b�m��Db.���V�Y�w:�`�մH������;"ƹ���Gq��S3��2!�����}��Wnj������q���]5ƈ�_4sp+����/Γ�o����ȑ���ԫtc�[���#���+� i��-B!׆sy����'�s\�C�ב�w�u?Z�5��S�q��i�hƃh�)Ģ�-��a[h�u�E�o���ӿM����i��Z���S:��nUhB��y�I��ď.��an��R�_{t��=�$�_
�W#S#��@��fNs���2�i��lZ4�mV�8��Xc;��nV!�#[H�Mr�ۦ�5o�;�����t�����uP|	�c�$#�H��v�dlN嶬�D�t.�e�<BOĂD ^my�vX���nr{#s�]����G��W�'S��}h�/4,e5T��Dh��H�hQ�8�9��i�� ��Uq(�UV�����B��=&���ҥ�]ٛ�j[+M����u H�q7(d�����6���s3]a��z[�j��^��4%�2��#ZB5z�br�%]�Z܊i"��^�X���aR	�}u3 ��B5fKcmI�J�N��E˗Y��!��u3crʉ$��A��Y��������jz�rćQ F@#��*�̰8ˍ"ҬYiO�u�m��'�ɷ���B9�O�И�\o6[<+It��؆T�/�bDڕ~Xx���6&DzZq��U$"��ܳ%�'�����ʆ�/I�r�<�9�޷z���*n6i�Q�d�[��6�͝�o���>t���`��Pbd:6t��)��XK0H�H��ɻ���|Oĸ��Y���"�$#IZ�"C"l&�%���� )G�ڢ5Th+mu���I���[F��{ӌ�h�J�%7�$�
������1֦ �G���X��F<$��)�(�H�?�@��Fca�!�!�-w �U8���3tnn�N�*|�b�8L�g�H�8�[��>����^Xt��}֎��s�����"_�V�Ni�pt:S1���9��fBF�i4?/�)� H ��KMq�K�L�Ľ�ؤ1�S3�ه�JJr�q�h�D)�t�0��.����ۣ������[N0�=J�+��p��O)	�y���d
|�8�����סb*4��l�+��$���C{T������Ď�s�ĳ1N谑 ��XQ(��ε�o9��P>ʸg�!�N볠,��y���9x�if{&H ��� ���tŝ�hK�%3:�Mlx���>ϲ.�[�V2k��u�k�[[�6�ȉ����|CMq4i���Wظ�7X/4(���������>tR��}#6�����t%X;Yr���%�rTк�*�AL������l����E�+g���q�vjB���C�*�'I]#�)rs���by��pqĮ<�ӁL��Z�s�P,�:w�����2G����y��8mfq�>n�����v�kGb��gfq�yك���y��n�ELDIn��}(��0�,�%�6��f�S��:{���$�?y�R��4=��x�Q�'ޙ���(=ב ���3�b�y��\q�B���wD�8���5��W��]��J���t�O��W=P����a���b�|�9�-
�b7sD ���I�l�@hܩ�F��r���w��l˹�s�
.�e�i�YС�ۍ�E�ܹ�S��\�}��+��3���@˴��]�@&�w��������!�r��]c6��XC��g�<��w"4?g��m+4�Tg3�L��穤{z���������l� ƶ�����ތ-ˬ��GV�I+4��˵+���3�;�R�! Fz����$����$G����gi\C��$#L����];�CI`��k���G�j�g�*}ef7��,�d������<6�s[���B�<`�@��[ƜV/8>�B��+}0ԶwdS������K�h
�E��L�L�HErK��}�@}��QJ�M3u�>���k޾2L3�[TU���ER�����à��
�dg���{( A:��L#~M�u���~�vHY�����o�4PT�c�u
���vr��F�� �l-g�}�^3���y���Q���xb.14�w�*6Y1��R�6X�,4>�6Q�Hͷ/���F����چG��}0�Xa��N1��I��Խ5H��׆�������t���e�l��Bf᱉|�<�a��pԴeJ�t����B;3*�S"�0DT�E��Y�:�p?�����i��MJm��[�塨�3�-�Ʊ�a�,�5Ku�i���j@,�J:V)p�3��D*[�Z���b�\ˠZ$2q�T�eJ+X��]\���3AH�����6�J���\��p
]c���rVf�%
��i�#���3=YCL�����U�1W3F莱��X��v��J�����0l�L^��Mm�r�������!oJN �wS�  �b* -U-�{���B�q6����5��[�\�5bF�+���K٥�(i�vg��X5��\�����|�߳r��A���g�XO�Y�8��{��{Z
�0���;�mq���r��g���!����]��3�_]�ϛ��/��8x~�9�z�g�2�4�_��5������m��Dz1A}y�x�&&9~�֛�U$�Q)��os|�ݟ��f�t6��>xu;�X;�+�x.w��{/`��w=	0�\�^��'�-<����ƶ�'�zzε���D��!�0cN�<�q�7�p��Y���K�=���OU��6ֆp(ԷDxO4Q|�usw��d�m|z^�>����k��-�;��M�7��oc�2|��*vm�>K��EŃ��nh�w�'Ϗ�U[I��f4}ﲫE���x������Q��9H�VT�%��Ď ��7b�j;�&qZ�s��+�&d����w���zO��7�]��µ���?Z��R���:�r��4B������pЧ���i�ɿ����˂̓;;�Y0�����"ux�Cf�z��M���sۗ�`D	f%R9���\b�ɴ�4��~��	���-Eh7�[{�������QDh��X(�Ztڞ��$��x���Y�=�7"��P��}ߍ�أ<�싺��W����xo���7�Ju&����R��"��Bu��1�(?}�L"�.].���N��g��'w���]�:Jf�M����{�Q�L҃�ZrR�3^�_B������ˤ3�}q��yܧwb�ݟ�8��#w��5����gkm6&�ѳY�w�������dF���!`����,}�io��=� �������l�n���yEI�8�ò��'��T5n�g^�L���kxV�؛���}�Uy� ���g�z�����i$_�����FI�w[3)1�3��sv�؄h���{!)�1��ܱfQ˪.��r�՞�'�xK����G�����K�ȋ^�H�h�
j��$x%���o�Qi���:��sݎK�m��S�%�$��V3�D̈ﾚ��=|��V���yV�^n~��F+�Z���5�oX����OX���^AE$dv�����+z�ϯn^KK�1.��7^�����ϲO�5[A.}e��1�>'3��_42��y@UPѴkVg�fc���ݯ�d;n�Gw"����Wo��L�?yЫ���$0�
�RB}rՉ<��𲬓����um�:�&׃�"�j+{��H�&f�f�Mt׺q��a�[3r���5�}��F�arac�ņ`J�@f�3�;^�ʣ'kO��-uR]��MC��RL<?}�8��yU���'H��1�2�W����h�P{&^��Z�x�g�܏�i�8@a8�p8�@�k}}��~:���m�e�
Cg,�Sk���[X�s��Ų2�GL-60ۨ�M��Д�����?��3a���I!TXT*�cZ�{Ȉ�^[b�U�f��1���B�!ƥ��wZ�I۫���r��r[z��vJ?0D&|�<��_2��x@t/cee�P��F���~�Z����/��/���|�����欜��~�3�0Lm�4�Ml��f�A�x��0d��D6(��_z�	䠼�Nȥ�Ωѩ�c���Y5��a�}��a�X�M�{�����:3Z�y뫻���uV�����4��E�������谐���SIx�K<������x٘�=ds���x��l/�ζ`И�լ��LF\�{���ۿ�!�
�A��o̤U`�Gv[��>�û�j�� ���3��1���(�����`���I��"Y4Q� 娰�٣�px�8Sx�c̼�/��ݛ
x"T����Ζb��l�I�n`�P(õ8D��~�Ͽ��m�F����
8\d��Eж�K��SB0R��ݬL�aJh�[uf(�s�.왘9��S�^29u���^&��%�:4Ј.������I���7è�$8��뷈��*��4oR�.&	ٓ3�,�q� %
ئ��tQ8����t=]���Ns�C-}����� f|O��t����̿���u���]��g?}�e�#.\�溑��Y���A�c�g^�,:�|#�ce3���X�G�,F� ���>hPV�BdH�i)�_�7���ч�>�ϻ%5\ku����Dku)x��4�0����L����5j���x���Ͽm���*ٙZ�z�cv��+T�\��g\���7Zk/�xP(���Xvӏca�����)�1ކ��)70��hD���va����7f0+�v�E��#f�2/++/ow�$������5:O�TES_B֑�������K�E8�*�����._���|�C��e\��4�H\	f`DVf.�0�ml�#D�)��^΀-([���ҵc�
���$d$[�VX̐L��V��Ft�Z�%�RݭBT(kA֔x�i�c��KQ3�HЙ\�ev�U�������Z1�.����M�+e]r�&"�v����MK	�J�If��6��
��Yt��p�)XkJ�4�u�0�̰P\�����WW�����m�Yx�L�5kKvSmiM�p#�-��$�
J����ͻ\K�]j�ݙVh����-��z ���`ـy������`t�4k7�:�c�����r.+T����8�I��!0r��N陒L��8a+Dq�\"_k{�^}�k]?ky��TAF�UQ��S^��Z��?����"~C�5�U�$�?Y�KK����%�v|?����(�5b�܈ d�(��" 3e���hB.�@�*�r#X:�"`6� �~��,��8n�Ǣ �.���dV!b��aD3��I�u��5>�'���G�
�������	>�f������C�GJ2�Sj�a	�2���F�ͩ|}��x�?��ק��}�&,�e�w$'�ttFF!�s7	���I�,	Uj\����Ҡy�6E���{e�/�����~�t�6�Y q�N�H�ڍ�TF�Af,�]Z���ћ\gu9�&�h݃L��&�p.a����F������-��h't�y�wC�0n���\�>(�<�*�@��d+��`��8JI
�����Ӱ�=V-��;-��UG�����+|F�5x��K��:�!�N?]���I�mk��Qr��L�����"1�H�Sn�CsewܘB�h<b0���|�!��k[w���Ċ�cB��E��c��5��U���?J��0�,�a�2�Z��6MWOd�da*�*U�x\hP���w�,:E��AZ�;9d31!G�; V�]hnP���&�l��KB���0�m'�??7zsB�ygr�_[����/�_��/b�7������}�%�"�Z�׫'��߼�;x@�ZR�F03�/Lp.�Q�5�:3
nR��X�;zu���2��O���}��P��YL��Z�Vl�oj\�j�ѭ��5�ЦLڴˑ��gwg[�z�@yS���0odp#bIn+Y�ë6zO:���u��H>T��mP>�ùC2wr�ݜ�*t����x��B�Olǉ�$�A�4���UXЄ�������p��CvJP�"50�fH��e�ԇ(�R?���׏u�;6{�fd�1lĻ#Np��6SxQF��i:!���m�\2T����=�QMw�8�R�i�]��((��K,����q8ʔ���5�K��w�sz����Z���4���mhU���q���B}+�<�iUhU���B���O�鉉y�=_h�6W�D>w%��� ɋ�K1.\H���H=;R�� �����)&/��!}˃�-
��N���`%�MXb���-�VQm#E����}%��ѓ��_~�潩5Bk��������=�p�����Dkc��\�hS�)Ym�(�@B�����m ���y_{�����o�ꉖ�˲�VX�L˙�K4eiJ,��s����spT�4ՙS	VpHp��zL�qb��*OZ�/�A�*:�.Zc��.7�����4lܡ��W��qh"����-�M�䁖���S��u����V`��PC׼w5&��TAH���	��{ݙY�N��~��'�fh�^�3�����F{ǅ_Ǻ��@ㄠĉ2LfI�>��X�wĉD�0F���xpq`)P(��JG��P"2�8�G��9���0���ai�IltK��C;�������1�/��\@E�J���N����f���ݭ&1/%<�|�ߴP����9�P9r����v/����u�K���ّ��qk侍�@$<G�>b�ҥ(#I�W��iih+�=�������5��7*���T�h���X,��Y4��bY�d��IC6�V���;�@���oG;�x���]n�MD l�"�f���b�F|��(���q�JR:1��:WZ�J�aF�V����B����7�j����q+�@s(˴�Ͽ��g�����	7���m���Hp��|�ģi`.l����=D9�L��3�{����	'�"o��"U�%bf&��~�k�l�k�_��
R�H�'"ll�<3܅Ͻ\_h�4�����0�"��)�p)-����֖�}Im;;L��ӈe�l�4�n��P��>> ��[
#���P�BΊ<��Pp�M�N��=�Q�Ԗ�w)�1t��N���#slvCnm�m���Ix���h�;�
�	 kw�Ν���2Z��Ko(O�2�f�L靑	�,��W/�U�x�A�����L/kJ`x+C0d�aS�'������/tsᘐ���Y_\F�񨺊k^/Ub�edVY�ۃ�s~3_d��Y&M��+5I齑Lĥ����'��~���A���ftS����۱�o���{Fn��#��U�=�&�]��U|�=�6�����o�w�V��F� L����S�ʮ᝻�L]���͐��c��[����=O;!�U>�|=�I{��m鹐�#%v��ٙ�.%n)�:{��Iҧtp����( X�%�u������dK�	^�D}�Qi�m^B�������h5w1�x�:� �?k��	�]��k�e,�yQ����U��.�Ո�<}�'�z���v-T����Z��l�/gna�A	H"Ҩ����L�2pd�U˫6K�޻ž��bo�m5�o�����^�n����b�W���V�(�y��v-��p�1,<9C�����#�_7�^n?=��6���H��~c$/�1fT�:�|��Y���J�Z�����/5y�"���MV���$WyvP2x�[�|�O�M��[�M�����x󚷳�-d�K�	���r`~�gޮ�����>�_(W{�#�ψgA��+�bp�ӄ�n��:E"4!�g��B���O_S2�G�@��-��m	�i�����B1�+MQJ@����%��8�j�3p����X�VҦ֚��6�I�bD#B��Z
�QN4(F��i�����-!�ܔi�-
�@ƨ��lh�F1���-c 4m ƬH�u�ެ�{�SE�(��m$�4�X��yqm�m��D*ҴЪ頍j����C��hjqۘ��j�(uKcF&����D�/��oU��E��bEk�����z����z�C��5<�0p�(Ҍ�~�B=�7��3UNB�TD�Qqb)D��eZe�>#C�bH0�v�Z��<XۻE)�C%0�m��0�Ѵ!���'n(�&G7�O=H+���u�Oe������{���*5�Y��P�іA��K'f�����m�S��o�M�A8�I�!�^~��k�Yܨ�o-d
t�V��,�����5�)��J�{U#ﴏ��V%��G�w��ɜ��﹪
�Y��iy��ݞ�������2e2U�%�n6�jWJb1�1P��f�SB�
rɵ�qi�ufU�%����m eM�h�c.ya����V�2��TҤN#6�@��	l�l¢�b�q!eK�UZ���Q6�m�P��1���X\Z�2�MK����rao+v�����%`6�6�	\ۜ���ef��@�ڍ*�cu+օ7<˄u0��1m��`�M��� [)�͙ei*#rux�mԈ�&B[o����6�̱T�����kB�9�6\B�B�5�,+���a��H�H�F���"V6spM*��4v�1k�9[(#U�e@�:�r�l�Rk1\ �5aeΔ͸�+f��T���l�껬���E�j$[6#�^��WF�f!DG.0&�CX�@�[l�r��)v�]�g-��1�`�نԳC&�,�`������Z1�(8AҰVWT�T�B���`���(��i��FЙcC�v��h�Հ�T�à�q�KL��CYR�umK�	Hd�v��V�`%��q��W��k
�	�:��JRW��2�[6��l4���JM�e�bPt���R7]h�))(3j�J\�j:�ƱMa�Ԙlz��A��ɥ�53%\#������V�I�vx8�	�YU��h����.	�]���R�����)�aV7`���\i��	��s�T�0�.6e�vln)cͱ�é�i���Ҭ��L�V�X��U��QkFː���F�ٌ�V��J�il�͡���y�#��N��%�L@��5�Uu8)kZV�ݰ8��:�R⭚8([��%К�2¬Z��۹�ELe�D9�A��c�� �W1�^v�ih:��rqv���.rۗ&���T��l��`#�Zj�î�X��Ùiv8��	le�e���SuZ�l-n�1�̲�̠Rq,p�%�+�Ѓ��-���HXcVTF��Z�Δ�QWb���A�!��ŵQ�H�\h�"iϛ�P,G�=��bS[#���a��j�����i|\5�H�&U񉿐�:�r��ǌ��P�Y�hn6�6�Dɱ7��^(Dec�ǒ7�<��_f#栥�n�����k'�����}�����W7dkڻ&��D��X{Y��VM1;1����G5�4׵v�֭[P�B������H��j��:��iM�q�H��HM��T�ْ�kʢD4P}�[?/�R$�d��Ӂ�'�Lwa�Z���"!�o��gdH�(�"��i���2c�Wo��^蜞���GP�k	���m��L�̄�|�c߯zx#��s�T�X�ɮ�1�
�cK���X��[Ai��ɜt�\����ZYI�j�nE�V���m�{�ae�!v�JVW0B�Z��IL�X鲘{4�[��Th��s��]&�c,HW��6^�d,,����a��C�i���0���՘�D�P�ic�Ųeų%w[��!��*��ū����%Յ�vXք,�"�ړ:�!���T�
K6�		^aG+Wⱊ� Pf3���-���Mæ��� 6J�� ��l���Եii�QZ��Ѳ@X.�Ciu�6����7Xf:���5m�+(�L�;B#���gj��7y����v�z<�CxL3��g�%A�
��}��������u<^������F"�J~!;|���c��3����������{y��_"^bh�6m��V��uJ8"�)�b4�eBg)��	Ks��	�gY�-SX���qL���0vv7�U~0�W�/�'�
�ӵ6%��i���^�4x#8�ʈ��B��4@��䥒`�E,��.ƫ�#��v�~��{��g�ci�oev�TЏ�ۙ(Y&��Қ����`^��O
��ۜp�~����q,�/z�}2�p���R���~,%�_�3;	�ZN�L5Te6��>>�W�{g�~���7㋜6h3C�^Z1���l��6���;��t!����X�H��XE�����������-[�mt�)/�H�ռ_�h�,��0{�4�XY@AZUQXĪJ��÷>}.�F�߉ Bǿ|��ۭ2��j��!�dO��}�u3�x�\�rx�j�B8�h���.��5<v�s�N�I$Ak�B"���<�'5����mL�8C���A ���4�v�܆@�Ӡ����O��;�o7'��f.ay��	2�m�5KE�D�����f�G�*W��YE��8H�r����O��Ӹ8Ӯ��镪�'t�b��v.�$�I��m5�NET��K�?f�C�\(x�=�Kwf|�>O�S�Y����|"9�?�^錔���څ�p��tx��js���<�!ld6F�b:�a���$��������GZ^g���h��>�%����_ߥ�oln��Z�t�Ab�ZV��C,l���zŕ���*�K�]x�����Y>#Y`4�rH0��q�$�t>0��#��Bݛ'�S4����x�����g��F�6�7�ϫo��p�`#���r6[��$����C����<�!�i�d<�-�Hmt��=\��C�'��k�`�9U�B<�#ѕ����چ3��a�����=��BATn%���ֆ�	�:�,�"t�����0r��-de���+#�"l�S�k~B���Q�>m,��p�'4���_K�&�{e�(5$F�H#sM�%�J������%25M
r'��5�k憚Z�����"�(�
I�wf�]͎&�9�~\FT'�)!��H���(�4/����+h-�TAj���4��kw�/=곷�ƶ�$=�,�&������@@�.	��4=�j,�;��옰t�H� �6�f%�V���P��摽᚜��� �5�$>�#�!:m��<�M���禇��Mm�>|5�}����mtv�m��Ȭ0��+\����LU���X�-Ո����*[.�c{���X��|�g���tz�ל����$G����C�m;�9B�Ƣ**#l�H��S��>��p=B�~A�*���m�$��B
�����C)}ߟ��}�|��=��m��tʢɯQ���Q�w�-��@���Ƨ���6(_=�6j��EK�RF�����>�i��>�g�G�df}���X^�RF�ڡ���#���@����7���q�'�r\V�^w,쓔�
����,��3~=ޯ;}(g��Y�-n2��H�;���0g��y���F%�q�W��\��l�N]{�gax�7G,.H�3�hN�j��Ǫzl��ջ�6Z�=�HR�-��dn�l4$3bU=��w���"2��.Sk(iA��#S,7���M�(b���er詵��O'�F�O!<�}�mm%�X���	�������&�@�5��	����	�Խ�'Շ��S�@���j��>"���Q7r�]S���̢ܺ�3��\�5|�̥�r��XR�u�F��i�F84ֽ�~���Y�����!�!��
���dCci�)��ޑQ�_is�y*hlm(�
=�"'~�������~p�W=���JHO�&Gl��8B�@<�Y�_Y���s�h��Ç��G���A�}�B���<��c#Af�sϔ����:�,go>��=���P�W+�O�za=������Yѕd��Ta!��e����o�{>'{��I�U�;%��N���{ �ޜO'�y��(-��M��R�Ȁ�����v�E��#��H�U�އ��%W�m, O}���c����F
~�ԳB|�D�=���z�8�s5�����I�}&�|��<Z= d� ��m�mĝ Щ���(f�?�82����W|�DH�hr�
#Bw��]�s�:�BB�#��^NW�����
X�uݚ��mCa�;�9�y35̀�e*+Z��`_R
���^W��;#�n\�3��q�6;*�4fn�ktp��lέ���I\D��
�5&���!�̐h�5f���t)��Lۥ����]�����4�hq��e�f,em,6(�\�˘�����i�#��eѕknClhٵ�^�2� �K�X\"���k�7�c�C*�ڸY�׳E�6/W8�1��QM.��8�.����[��[%��^����c?�R���.��dn뱼�h���b��ٙW;3X��*9t����+q[�A�[D:�L�3&Ż���} w�r�Ĉr_�"U(4k��M	�ݐϜ����7��SH�%ED�����(�!���ac==E.���������2��˹����z�ɾC��u�w�g��V�>��͡�y6t�=�X���a}�#3�}��g�9�=ooz�??���b悮�S=��f�@�ͳ<���q	�������U�����%Y�f��F��Y���9���KTh��-
P�|��2��d��3�S�L�!B���8Gsl�~|�l�έ���2���M�w����D��w(J��DHBAH���{����4�<���]A���W(���ADf����SΏ�}Z	����B���K��-H�=���:�(g}63=�J��]�:_&��(��J��$[�h�����,r�)�LU6�-H�p�ah�$f�iu.B&����Z���[���6?'�O�iz��(�5�C`��a*�G%�+e38��X!<�~��}dU�Bȑ$0���}7c����gޅ���·��,����1�߉�!��?i��h#a��V��ȩ�|������^J��նL�K^�m�|� �S�J�^٥'k�w%�q��H��yTPn$�V7�� _�rNY����0M&���w�@F����i�g���xÛ���E5끺"L�<���`#i�W��;�GM��v�D��g���:���@�_�iMk��gq`a
Y�r�)�Q����Pe��%Y�}��K6������#%���-��I��I)�Ŷ�<g ,q�8�P�2�Ha�ޢ��-�Fi�����Hh,8TzA'���8������L�����v�Uݹ%�*(������,:vx8��B�*����:/��gFP+���\b�YHQ(�w}�,�(Ly���C�A*("Y*���-�.��\-����,�.mu�����F�miw=��BJ�X���0��V�\>>M{�͕�Q�x�5z�N���}��x����wq3����LƁ��8 s��w$�h�
���}.�u*��g.K4:D2U�������^��+ct ��u��Ę�}��9
��97�Oc�Vu��(�տ�pe =z����D��Y�o0wL��^�d�6�\h2j��'�Fo_n�S�N�ܞ^N'�gM.����C�/v臝gNi�t�����8l���l4�R��Q)�v�e�_���Tx���ST��-U5�+�v�;F[h��Q[Ҋ*H�Pi;
��䗀H��i�XZʴ��g�M���Ob%���r �?����L����2�Y@A�X��6�x�CF��35��'^�<�XeF���	��'�(����Ձ���a���#�!�`��#��8V�O�@@!��`"]�OYZ����>�+��@�Cl���>���	3�>}#f�Z��tX�X V�q��q�YG14�tQ�.�ЎC5�l�G@��L�2cra���ĥ��K ��QL��g�w���`�v*�J/~(�9��8k�O?�fN��]{f ��J(��$(�þ��wp���7�e]�]�X�1�w)C��0�}�|��?��)k�����L�d9�X��4U�|�/1�;��Y��͉_]�톚�����u%�uj�S�%h�f`C����H|8�!��� 1�*�6*�k
;41<�<��5�C�0�Ӽ�<;x�>������.Ic%���i�8��S��~0:Z���}#�H�������i�|	q�c�V��֊6l���e�&�!S1OX��e��4*�b#)�Y�]:.���6^���s�I�2#^�i�����߳}�����i�4�,HҋGP�K@�%x���㟿X�6?{�3�?]�-32[�wZ������͹j�`�$����S�MW���EՐcp�� ɢ�~��@��ް҂����8~K���((����t~p����u�����5�,1�5�v�݁K�[����Y�@3vV�?��~Y��.)�;�BJ��f`�(K��P!d��<SF)@fAͶm�G-S���#X~�_�ˌ�L�f7w,���U��x�,y�}�-�[�:x�OX�x��p0��gVĉn����OxxFnv��>�{��oݎ�q!M�F�t���&�E���n�� ���*G�U�{���UDF������bu�x,�JY�ܻ�d�ٜ�`���"���08j����J�v�9��H�(hEg����{ts�I$d���fg�BҥC�Iv]�0��P���}�c�s���;��E׮=9�<w�Ě��:V���'��W՛*�꺨4�UDT����9��:ZG^;��	��.�ٖ�f�y��L��/%��#\]U�����횷�WsY�����R��C�|��	.Y�����.%�F6@��@)K��X;9A�1�T�UJ�[��˅���4h6Q���L�mc1M4ee�:�Y�!TĘe�\村W&���ui�S-aB���F�.�cBj�Z�d�BEw����s	b�] +G���;c��6�12���t3�նذ�%�X�����a��+�g�oW$�m܎��5Ns�,&�V�PM���Z����ƚ�K"
�JC���_��Fmt"m��m�q�����R�I�K�����v*R+mce�k3�r�ٰJǋ%if*]Ժ8��!�1s��3�
����u�^�`�"4�7F�������T��N�L�l�tk�z�g����p7�
^x�RY ��g�y$�Ovty�k�z��a����pGZ]1L�3�"�0�;��������"��MR�ԍ^��τ�r�9���r�73<�cy�U�G�U��gq1!��:����\uEGdn��X���,��u�H'Ī��sR1�9�nU�zHT�4�y��&��%���]@l�s#�e�9�c�;9p�Y�'uwn���q�$�E��=��q��9Sd+҃1��!����H�d���+���4��Q�S�Z��_���npq���Μ�]�X�#B�G����S#T-���6Z�q#�d8�G��#������ԁ�Ra�η0ָ��ng�`w�=��̣L��yY���:�p��]��z�8���ʁ;-�>�f���4a'?%�~��i�!�:��	<�,���Z�X�㑰-'�º��w�SX5��Ʋ�g�]�{�oE��^��;Y�������!�~A%1������� �J	���
��;əQV��@�S䍥s?Х ��W����F��}}O� �G�O���'R������O��qh�c^ܒk�n�F񗄒M�)��Ш^���j����f9��Z�W8�ݷf�H�kA��P�#��	Ӻ��Ɨe�'g!ܪ'��M�4T�3�=S�~.���6�� @�����zqr�ku�XM��b//aHQj��:�{�I��B�|���gv"���T�=(����`A�� �K�T��;�ox��10��j4�g��`\��/^	* H)%����8��ݪ���Q �L�Ee��[��@\�6֣��%��m���;rd::�ⷈm,t�gW{4�]� a%�{�@LOp��=���z�2�	tH�~����߾�?��u0�-3-h< U��pF��ʣ�U�2� ك{���*9��1	;��C4� �<���Jv����;��<n�\�g%��	�\lTe��p�~��~���	�����pr�7m�ߣ+zD3z9��|���[���TLQ���{��á;��Lrh^��l���׽��?iZ"ܩc�-�fW��v�9Ek�:b��1���{�5��秣V�?Y�{�[sWc�7�O.�-��{n<FòDw%�n0��%??m	1��?!�6�_���%�zjb�}���>����<�5p�2a�������N�5�'f��l���L��(�|��M$BZ^���m���}�=w=�f�ؓgM�
�)�6�E����0n�e�Kf ���6%x��f:֒� �״�nt�L��*T��v�;2b�4�@�>�zo=V]i����'܏s���>g����D��W�{�����32��a�3vC!1�m�off�k�Nǯ�x��XBloy��f�KM�� ���j�ܪ{���zB��Q�I\��1,�ۍH�����?�wwX#?�jv����j�ۈ��s$y�����k�A�І���26~(<��˭�+���`G���e��y��]�|Vr��d�7?w[��cܽ�� ��nNva���9�v}���sQ�*a��6'�g�3�e#��oXy�8!��1�m��7�Y�������Ǫ�#�A�
�ϱ0v	���'g���a�u{��~�b�;�=�}�i>p�V�	������A�����z6~��q��]�]�����q&�L��Ԟ��<��	��8v�����SN�?!贸���f+i�!�XG}4����	�������SvM�+Z��m0���Pa��i���.T:n�R��*
z�ұ�>��%r������E�Ĉ)��AEMzX���!��j\���Y��ɩG�w*vQP��G!*=�m�a+$5�����Ĺˢ[6�T�7�=%oN�2Q��_w/|��V�32�d�w ��k�I�E����M�-rAc��(`�j4�#�C��|��X��0�M�RW˩V�)ƌj�����̾���N�����\	�Grvz��\�K���LV5���*��uZ�z �M7KGw-��*�QE^�m��!�R�-c�D\bR>bn�׬-Z�Go>�+�F��}5���B��
Níܪ�Dd����X���h�H�B!m�b-m�{�hU[z֮o����7�g$hlM��KY�I�u���j�_K�+���%����[z��<���[�f����"m����M,N��QhZj���������z����+u�b������� Y�L��W`}�a��������N�m��d�
$VFh��z��LxxJ�î�s9g.Yܠ���~|�,�m�n"��\�AiT*$P{^�����&�P�
�9�7�߲�4MEk�-n�l�Z�zKL���U�g
[����m"L\�[XB䩶�cir�e��H��I�~ݼ��lJ��)�N���z���濺U��Ci�J��w���W���a�Fˋ~��%kr(;:%�Q����q��a��G�r�J[�-�3��z�Y��r#y�����4�24�\.Ė%0�{ Ȣ�7G^�g@�f�c����<)��zR!��6�|�����r˻*�u/����	��%�}��wkgM��]ڮDˑ�'����+P^�8�"��r����<K�����r��I�7�p��)BV�x��ΐE�k=��o�}��f�����45{�{�'�{��4z��1��	�DH���o��k��e�k�f;7dex{�������X��M2֔�V�m�f��vt��1�A��L�^-�.+ �kI��(y���ЗUW%ٲ�����d��z��U��c �<}�W��B���6�O-�un������'3�S;�;2�^g�N�t�t�f�4_��̨t���$�������,K�w4T�P7+D��L��� ��BN��d��y�F�*���-F���>$B��alԩ��IVB�����7��8ۍC#���6T������a��U����)Ͱ��}#��_r�<s翳����}f=�o�[�%��zg��I��X��H҉�b*v�ڡl����E�٫��zQZU���ϵeUH�m�Tֆq���uC�R��O=[A��,Ԟ�$�0s1�R�c,^�Id���T�}��8���zv[ϵ7۷����[x	�%\`-,!��햂��"*��H^�����|;���|=��u�!�����m(��e����S:����f�
*��!f�xaii���T��Mkslk��	5M&`.��G��%֤���Šk-M���0���]��!(��6��m �mM!J���v�6�%0�%%�A4�%@�	\ �ZX!3y��\�pC!��XknW\:e�r�#�n��Ћ��j0�0.7]*	GgK`P�B2�`%��т�ғ.4�M��r\�&�EТ�P���!�٦,5u��1X恷j�M�ֹ�n_�7��{��-D�+�{��	m��wDW_�;�gz�v��)�3�r��"S�󻡣 zڍ���Z�EBr�>qO�,��A��5�J� %CD����L������I��J��HE2g��/�u��e�T%��ȼ;�c�c[�T9�q�C�Sg��`+�=����a�X��O����w	�s��2�uA<�OXv4l�W������A����lHp�����M���bhLy��kflձ3��6	�ܧ=^o�r��;��Zp+a���_T�;�^e�)�fr�`�u�����e��l�ikf�қ=�+��Sm��lX�m6���k���~�׹�������)j��Q�f�R�r�@�G���<�wl�� �j��Y�fw`��v�&��2;�j�m�3��LϹA���-���f�zxgn�T��M�����'�N�����z�%�zN�~_�79p�L�"���}	[��[�q�6P���n�"Е�kU��xD Ӽ�]�,����oq6[�g]��f,�;�v,����v���.�kO��`�!�C_!3vT��}H�SG����t���=�#.�m�̻CR���:���,������=��v�/z�g��T�쾝��3��i�6���6�m}�oܓk��u#���]J2w>L	Eٹ�T���\؇��	��40���[`CT�1�%�e�D_E9Y�t}L�a��-ɒڰ�hK(����ai��5݀�m�h��\��Cb�nʓ8�q�]�H�Nc�XJ9�J����h�k47��n��͠F��w$;9tΓ�r����Y҄�&��v���"&G��I�@��r����}>\5SF�u��uٸ���-zs�(��D��8g</��q�vX�C&�]��fb�gv�!Mg�#�x�HCW6�p�n�	�z׸�cvj��V-ݙ��v=]9���2��y�yN�x�d�;��O�}��}Ǟ���\����¬Ν�YDc�-�P#;:���-��'�W׸BϜ��d)5��2¬�����2�9�߮I7Z�%�V�:�K��\��P�jDN5��;o��K@�1��D0���X̝����qjY�&fvJݦ�8�F�1S�Z�UR����n���{^@4��E��r	�|~\�L�L����vS�qw�HV���S2E�o"w)�,���!�.�Œ����[�_|d�x:�C}Q4f]�oa�jې6�Íq��;K�G�C(�jr�]��Ȕ
vM�y���O���ﭚ�﨧�᧏����cOs5Uڵ�M[�ZGtk�فsg&d�p��]�ãB�}�ʒek�������35H���1W��_ڒݹV
��:N�s�1��M��l��Q��(�T]�Y�o0��w����5J�J���P#$�N�U]�Z-����KK�-��D�N�F��JZ)]�*�xV�#��ڮb��t�c�왟��3��Cp��ZS��(>���}��L�復�K�nVܾw
 9
��vM�N�����A����:�q�Z �A%�Za���<�`��VV�Ge��̓�ᅘ�O�,l\��R!��$H��?
����>��Z�}�l�=�H�q6�Q����B�~�>�G�xw
7o�����P]����\�t��l�zR�F}�C,�+ڎA3bt��p�j����˅6
|Ŭ��ݻʆ�T�=�4(:�׫���}�$n���Ӓ����,刽m���ak����b�k��ѻ ��Ŧ�)
:��y�{u?0j� #@��N�ISޮ����N����&d���_@ޡ�YI,c���=�ʅ�6㎦Z�h�a��@��\+��R����9���*�*�֪��WV�]��@�S�>�0����ݿ��{��~�����{�ޏ���%��Mm�U����-��nY�-ĥ5e
��L���\Q�0L6�u�x�cl�93�䂘t�cͥ���
]�Z�j�5��L�I���v��ʹ�n�%Dy�R �%4�a��� ,�� ��4e��]���u�Ы�R�:�Uvi)uz�4�QbZq*��
�b�BQ��L�څ�m����sf����nt��PM�w�My7�s4s\!�����P��@�LR.,U�4͵1M�ͦ��#e�i���3����c�{O��Г�I����)��o�q4޿K�s�K���������I��O�����I�T���@�7bk�DU�Lox�=��Z��6�o��C�z�f�L�3�����'b��t�ֳ�Ŀ��,#q`����Fړ:Xk���A�̝�9gfft��b6w:�H�4gM�
���M�}�
�v�����m�}�}�"4-#Ts��{�����r��!/#�;��/9zD��k���q!���?b�\�F�T�N�����Ù5zM>|����X�Z��/m�we۳1�!�m��6X�BV����֚ڬȍ]0�%�m
�b� �sw���b� Mm�Ԉ����;�2ǱÁQA�������̻$\ؙ�}g�����>�&�.U�wmj9�v����̺-y �VI+b�e��k�|d�l��i��Ӆ[�E<��1$�%\��QZ����:���} ��zŋ	�^vO�WdM��ͣ��*3��*T�"�N�d��+���.����i��E��"��b�[̽zz�:q�w�k2�R,Ν�۝��gK>��Or?��pNhnF����w�z��v�҃J���KiԶ��㭞۟I
�eDظ#]���{w˿b}����k���?f������i�u�#T6�O��u��r�����ē�uv&-�̎kZY����8E�?��8�3E�ķA������[M��ˇ���*�v6mc�[�T������}!�yv��Gk\6cj��Dm[�=E�#���:k:RN�~�Ϗ�}XgU�]ˢZ�&h�lX�C���Xh����T+ͧ"rEē���1�k��	�IԶݒt�3��f#�Ct^w
��bN�ne.��C�،)���ǐ�G䚻���(fE'?f1��߮y��J�О�T�DiE�9M�[9�Ģ No�DIG�G��K���?�>�>���$��BT����Sm��r%~vO߿=��p�Ƒ�(��x�k�IK{�K�z��w"g	�onh#rO���]��v%3z�C���9�ؓ��ߨ!�w���~O��{N��w^T����@�jC�X�V��l�\2�$�4m�4�⮰D���7����&�51�j@G%��>�'�%��O�/�g�5�>�*��X���I�x:��= >��`�;�b���c��Q}��й�����KE��m�b����v����q2 r��$���'�BvwM�;]�8�����\	+4�jܥ���*R��۷C85�nE	�"��{���U�_�Oď�$	�Keo�S!4^dGu=E�s҇�%!�9�vf����� d8�ʬ�#>�6Ն��6��U�2��=�)��m^n�	��kSM�줟Ø��o_B����[�)��Z���=������C<��P�i/��}� [�CT<���Z7B�k1Rm�3��70�j�`쓄�͐��r�\��c���Mb�����VR�eW�Insk�B����^����J~��r�p�N=;#�^�#�Я(-4�C@�̒���wt���Ç%s��óa��K����+�c\@�9O�f��ڿ��}����#���eq7���5�}s���M�
�ۻ���K�����'忡SZh��?Y�R��j���x��}���v�R �P��E O�M9aH���:��F�7��:�v&�DP�����
�LS�&I�tt<�y��b�g-����P*��i�d�;DJ�gd�&��w���/����F޻��_o����������������}n2in{�p7��g�~N�s(��u~M��[��y��pC�ʧ���8"�6[�fi᛽��$,󖵾�3L���r����%=��g��W�c���t�n�&qp�н�,�{P��=nwI�'V���78���rl^}W������{}���{}��&���97��&�}x��	ͺiN�8�zi���z5�^�H����O9Ybo{���w�
��k�3�b-�Z|�;�S�%��xy�7�.�{Z̐hUҭc��i��k|t��ov<Cڳ٢�2]�x|��%׹��/v*������ڻ���ž��ن�07�4Ag�����c=��C;�YS>1Y�{�>���f_?D�Y�����f��$�
iÙ�܆��2�羊��yz�j��K�9ݓ�Y��9�ⷥ�Q�ćh�{ծs5ř�gn����v����_�S=[���Ʀ���o�~����7�Dü�[��&11o�����^T��G��^l��[P�i�|n��5�{��af8�f�����{l��L�nvռ��$����#����F�%�Ͻ����������ZVs�\�pn�i�=7�m����e�B��%M
Wz�(U:�_cs�n�(��ǂ���Ozl#φ�h=�Q4����[�m|��`k[ys��^�Z��k �]���n7��tNG���{ۺ^�β�8�K�O��M�ƻ6ܣ��u_w�Wo?{;������ɓ�L��'�,�sʊ�Ɓ/�A�6h�C��=FEYS�,��&�8��G}���=N
�]y�]!c*��ث.��Nc������n\X~���؆	ݴ{�_�s9���"<�����k��o�L���:W>�ᖂ���5Gu]�Ƭ�c,]*�¦ř�D��:k���LK��Q�rh�AtM�����ܥ���:	�XD��ͪ�PY5]�wi���d� ]D���9"���[2Z��,�1�l�Q��%�!q
���u�����e�ٶ+��Rī
k�c����uE�õ��R��v�-���P�i����X,��suR`c��ِ��h�歕��j75e��T��%�V�%�m���V���j�rۢ�� �����l![��a]pD�į1���k�Уa�Ytcҭ��ظ�
�1؃^]f�֭P�fX�WL2��3��֡�	�F�J�m.����p�<-u���d]ƨXh6��k.�
��X�Sm�U�\�E�ke��P�ȶ\�k�h�l�K1K-l,q�R�E���D���&%�cG$���8�f�c�.��1-�	�lGK�R���6�j�Ժ��e��T�3B�Hʌ��k�c���6렶+B�d�)-�ˬ������սK\K o"ާ����qcYqn(����R֥`�0���[QKr�P6cA���Wl]f@�Ml\�m.�l6fЈ��sabFiVQ@�����1)�	��n��Q4SM+ B6
�bZf�갖�e��-�����)��T"�d���6�Mn��T�&��`5ku�Ќ�;1&���38�"]��T�:Ť��kټf�RP2��ls�0D�E�n4sj���]�XA�����l�WL1�wcb�U�k��\��%��5j���-	�Ƚ�Gl���,��mn\��*m.�@�@-f�еK�	enx�ږ*,Ύ�`f�5��C,iڼ�#�[�L�f�K�||R�|Im--���KM%�+ɳ��).hgh
e�F�5��$%Z�rvc���w<\J�'�ג�B,50Ab�1-�#4Έ亚Xv+�ve�Ɂ+6��vj&n�\v��3�1�SZB�"�!�K���c��]�`3���).�LY��%|�iQ>J�Z	JD�i?���7)j��"�q#�"���T䈭4�":����뵡i�>�YkP�i��G5f�^|Թit���\Bд�#\Ւ��1����;��։d�ݥ��5 Ҫ5��Q�	KM5r[�hw**4�Ҫ.$j�D��X���PiZU96��I�ě�C'R��J܈�:Y�Uƍ(���d��-�syu�Ԑ��Dq��3�9�$ ���i+���TDT�݄	"jTU�X٩�I������Т4,B �����r"�TW�����aPܨ�4"RV�@y��3!6������rcAfns�S��f8���U�\�Z�SVCI�iZi�CJ�i�3+���"#�ՐZB�4+���N�V䐕�9�\n���A��[�Z��k]���B��D$lL�F�|�kdRҪP�yw���憔���<$�r��HjA���g덀A��l��PDӅ�u&��>c�5�j�-���\�3i�YM,^��l��Ɛ�S�SV�k5Ԛ���̐��&l׶q�[����MHa2j��bnh�]h�%%�.+W���IhD�4u�+�%�M�఩n�DZ��.�6k"�l-��V���s���:]�mΊ�+��3rҲ�X�1�BlTԹ�.���$�5��)�0���("�2-��H@ChģA���0=X��p��"j{���l�ƶ�Kf��-f�Q���J��G9҆6n��=A�^�]�P�&+�Nmчkg.ܜ���9����u�ؐn������fL���G��.;EوM��?&h�Ei��G�U�Є�ŋ��-�#�f��L�:��+���E�JDX�\�xx��<�%�&��D��{���d�u��'S��h��}��a�]�.7��wh�z�wm�6)"��=�2�=y���U�Z䗌DW,��k���r����|2��C+32�q��h85JH[�I����fn�i
C�i;W21��6�C;T���!6q�.�fwG�ɬ�3G[Cs�ё��h����[uU�
��`qL��E q�܆_*=(��u��>2!~r(Z�N�,P��Z���w)����H�L����~��{ߗ��������1��xr��s)�(��u�>/� �=�A}*��Ү��9�yo"�J�������w����q<H�W�$���ې���_���O���w\4Ylf'�aI�nu�UL����oO�U8�6�cJ2$}뿝M�}�ۿ�ޙ��hj�'������nޑε��{��S�s�r��N_73=0���x�v�Cp>��q8K���=T�7��Ι��)�p]2�����,������Ơ��ߧ)��;�(6��m���]ge�t�֫�1�Z�11�K��k�m��.�ua���4F
볭m�H6�#6iX�n��g�~�#�����aѝE��43�4���S0�Hs�!�U���.��!&	�$K�\d��:�j�5���)�p�����������0e�Bg)�t��yؖL)ᛗo�wP�<0��+�,��iw��J�{�Vy.���ev/R���7��{�8�P����e�l��G��^�#L�o��S��M�fˉ�(6M��m&�����N�|�ė�)N噼]�LK$��XIaUI�P�m�W�5ᱢ�DB���4$ت0��yY��,Rr��:H���2��޼�#f㚝�8�|��qj�NѕԦn&H�0CϡWWj1]j�Y�vլ�X�9�I��%�nX	\cYL$��R��;L�]e�\��4?�J�ؐ��u���3]���M��1W�^�DK���n�lm	e��QWup���r����/���(��]�wyf�>¸�,-��ksn���*"�;_���`殘�`��e�����>к޵R����{�p�,,M��PiS%
�V��5��ψO���wS��mD�і H�)���-mH��s5a�3p��e\��@%�0�ʧ��mZ�kUw�'!�	Vj�<�^}3wt�7^�K�^�g��}h���>�$I���A]����ƚm��ӇMZ]��r�#`y/wӕ.�Yxg����㫺e�b.ë��0�S+���a�ٛN��ǻ����2�P�!��v4�A��V�<�Ҥ�[e6�퇜	���h	���Ґ�ٙm5�M�����l0�����
�0���
sC�l���ϛ�&0��3�0d��/��V�SB&`�A��%sZ�U��yw�B�d4l@"F�*�ٚq6I(�;X��4`���;��WJ}L�Ӵ�R��nᯙn����F}�֌�F�L���2�.�����������o���kߜ�iks蝃�/V�Gd$˃���N	LC�0�bcۼ��Q1�"�GC�"�\�Kň��âP�I>$	AA�҉��wܗS�%�a�R"�xT]���L�[1�/��iA�6[a�&������%)�x��AU>��ZV�Zh1gy��r[�.Iyh1.�B��W��H�[�\&T)�˴��nP�CDYmK��P�q��Ր�s�lh˷9p�\�acp".��6\�]�`�{2��b^�	��b�	���E�Mr��6۫�&�WXڣ�u4 ������:���b���s����e��R�����+.��;4�MF&%���l�4P��խd�^`\w�=���SFz����d�S�3��5��	{*ғV�����@&�=�	���ZsD�[�l������_l�8ˍao�6���ѡ�a&Ǡ���&T�(h���?O�����	��__3�q�bpg;�I-b�w�e�.au�kwL��rJ.��.��pk���^�\���lCF����:Ë(�R
-%
��)S���i���x�1����!�bF�PpB�a���8;1F�Cp�%hņzD�Q�$ O�F��u�k�!Ul����G��9,���lܯE�-:Uz{!�+�T��Ϳ.J��6��͏��>���Ȁr���A�z�&d
b�΃��e]�[�J ��!��Pqs���,lsi3��GGC a#�6�l��-��_��;7��	�)����Cx��ۂ_��y/o?��#!�P6���M�5�VW��^�0�{ɑgg�N�PeQl,�=m������R���n�;C=߶WFci����!K��6G����U��"����Zx\z�,��u�p�CH7O�r�Зhl��;�>���o��;��׻��9^��uw����:o�y�֒�d!������jbċ���q�r¸�t��v@�D�۾�c{��~*D1�h�$���3�����OY"�"��nF�ZwgD:gbC0(�=l^�4��cY���(�AкUu�r��s���|<i��z��Ϋ��.t߳���Yg�c��jK���bF!f�̶�a����6;�6�Bm�!V��b�9��Z�����t��d�0�T`������ł28������5�Q�(�, ���P���Yƅs��"8�]��������]C��}s/����H����1�V�D���x���.cxe�ŏ��?J��:G�:��̛;.��&f�:�q�G��&��>���ݓ,ѳ��7�甿i��/}/�}!��ޛ7΢
��0H��rE�W�ޙF�p�mK�y��� n��m���}����.���َ��md���L�����q^0��W��6���_��|h��V�{�|7z'��`���L�]��2,坜3��3�k�[\�Y�ש��g�zM���
�5��O&��3h9{�w�l.�Hft�(�L`�u���-`f3P�]2�.Ѹ����0�f\�Qqp̚�W�_'��O�{�y}0�������wVX%宏�Iu����Z{����,��߿�l�V��Y���3�*�p�J���w��,U�ʫw���݉͟������h��UE���꿒�*(�o�]��^G3'O��~�1�*��[�avٱX&(9:�X�����a�I}�wNJw)��Ddi�%�����g���\�g� ���|�.#Nk嵱��GNgxẇ�ۃ�b�]Y{��z��s˦��ff�=��:&L:�z��2�oK�fMM'�-S�o��s��$���ک`<G�¿E��:�ZCo�O^>������
3�ץ�ֽ�=�`0ŰbwB�=�V.B��2jjkl�6[��t�Æ8�2&`�
���pciEr֙�D��[c�bj4�n�R�pnع 2�~��|����M��%\���K$n�w��� U�b¬TB{�Ԙk�ɋ8wfL��&�����F��*.y�:Q�q5j�wh|��[��ٯ��y�JR�DE�EDE�U)E�Jb%RR�I���x�቗�*���g����7@iW5c_ED��0����^c��M� !ċE�����@��u#y��ˊSmN�����{D��j9���Z���h�p,c{ɠ�p��d�UeK��GL��zQ�j!�3���;�e�7^�⟆�f�HSzA�EC�1��1Qd#v�����#g�v�����t=�ҲK�`6��A��c�a H��%V}e���#O$T�v0,�˩���ZQMB��ȝ�����9�aC&óa\�b:TMtj�J��t]Z)@Q��YCG���\+�q	]�L���&�H�4a.Xm)�6Ո�Kya��4��!�JZ�p7\ʪ;d��a%��A�̡mH�jP����He�a�qc��L���m�s)��̶g9��s,B�YM1�CL&��$e���t�K�S'��W�G]6�����1�k1k�­V�쪩��-����f\�m�2˵�%�Vi��b0Ĺsqt9)����r񖅙���.h�ڱ���M�o����M�`S��l�b#��5v�!Ϯ�Ɔ��_z�F�I�2.� Y&Z3\wq��H���2L���[�я��s�y�3օύ}�}��5��6�M�~��vk�y\�F�C"RO������F�}'Z1��S�*���o��Џ����{����R��#m���;�@��ޡ�J��!�8P+�ch{��eANX��-�e[�kѝ �M!��:&r�a�#��O��w;��n�$1�I�ۯ�d�,lO��t�*���}���ʉ.e��j�Z��n�R�6��HA��W�l�4��j��4>�K畕�)��g�^�Xd�����>�xP�ۉ	gp�@�ʿ�Ȗ���/^B�;��軐Ģ�ᅛ����z�e�ۦ��3ܳ���X��>Ǿ�p�j���%�j�t�M����ɠDh�bG9��B���WA�1�B#��2ژ{]��g{��J�{���I�Z �����3=�����_�S����64|d6���>^��:�M��37�����-Ś.c���3����F}��24h��ǻs�d�Z"�fc��k DLooZJ�33�N�v	�8:p:�Y��X^PJ�k_]��\�F�:]�?�����*������*
h9;��hM��^�u�|������'���*�9�����Ł�]g<��q�j�[1Q(������F6baCl&�Q1q�%�L�T�~�|���5���@ZûJu��VpW8{!����H�� aDh��-�u��m�ir�Ɣ�����^���k���A�U����`�M��CA�AῺ�ϳ-Z:'�y8tK{�cC�2��\3�d�c���3�xuD��f�3�����ѳ��&�w���p�Y����Ƨ�{Vf�<��̷G�r�/���ފZ���i������o�!�8{_����ʼ���/f
��n�y�>��8��j��Ex�a'�}�ۓV�o{y���z�b�~�x��[���MT�;��]�Tц��V`K�>j�2^t�є�����8��Y]���dp��^��޸=�p�~α�8���1���fw�nv����ڴ�� Ł����7w�˱7²���O����������_���:��+�z�N�k$b���;�2q�8r{̭J���nNΣ���va �,H�Y��A��9�����cuG��LQ��e��͙��=�o��ݾ'�{�1sLI��`+ϛ[<�������4k�2{H��Ͽzn�Q��qvxXm�u��y�W�ͼw-��|ĔZ�����o���)]�pz��v��=�'f�o3fn�s<$P�^�9yG���Ѽ�&��W��[��$=]Ǡ�kfH:�L����T�37
dv�R���L�e����{-�"�%_��*f�	gj1	��t@��Id	U��i����p:�se$rÆ"I�c}�ܶB����7�G�5�7)��۷�t���}�k��J�>YTi4/��U������i
Q!*�;��]O�9����*���� ��+ڹ$Fx��#�=�x�=3Ìy�������R��<������wMw2Y���{+��,c�%mtzbD<s���FÚJ���oe�i
Ɉ�C"��qq&�xx����(��|̆8W��{�e�_lkl���?������,N�̳�Jn����F�I��il��Wp��0�+>j�gώ����- ���lm[�z����nc�L"n�&y��ߗ�$AK
~#� �G�4V>�̪H���C+�ac֠ڦ�D.���sQTÑ� �(�� x��kWk\�l���B=ʽ��DZ�1���Ϳ���
�j�����I��"BQ�H
�:Q䎕����Rh6LD`�e��X�Hvo�X�:J/�G�!P�4�F"��:�
��8�u�Y�i���]Ù)��߹jn��c6��.NX��	\���C�xD��KC�����O�!E>��aE�i3�҃?~i�	�!�lG��-�&'����߆3g�K1	��|��=�᫯�.��;�t��;�fZ&�>�7*X����9��(����S)�mH�+�=$���
>$�##d��ػ5%R?��|������B�@����4�D���_	�/�]
����w��G�i��H��f�V�Ƅ��gJkf�f�L��T#f�&WL�Y�[iU�k8.ȅ��>^ =�u"��JpKi�b;c]2k���jBL���4��X���SIK�E؆`���4p��y����pT��h�S�S0EU����4"0�r)�v+�c]x�����
:��Ļ�d���z�U)w�u��p�Tvyv�14�"��\���uY��Ml��t3K�0N��ⓒ��m�7��~�\w�����%lt%��+y	Er~�m;�0��^;���Ȱ�s �d��z�5�V��F�dz�QU8�R��9��RO������V4�R��c뼞�� m*"7D)B�O�v%?�:Q��@�:;��Bf��h�~p���^�2k}m���>��������}.��T���PT��Y��ku��a����^T��\��M1��v�c��1N����fu������24j�U��L'��0���	���˝�g�,�ջW/~��h�}�;��gP������^5F (�HD�T�ߎ~;h�|)c���e�a�	�[P��3P�ZUOE��:.��b�L�q�vo#m6�̏�:�]ۏ ��C�VNh�����~����7	�.����n���8ݑR:	���}:��ǹ�o�ɐ	 ����A�^��0mtS��p�$ݟ��1��as ���3�3x�8r ���G/Y����s���~���l�O��g�9C�]��<E*dQ�v*譄����a��7,d��dH��sv�U�����U�<������5��}ϵk٦K��ZZ�qb Wq�\ԗ1S��Yf�-ɓ)��Z��YX1L�{�k��1��.��IV5N"��3n��RH;Q��s���<͵�JrZ@Kp��D2D��A�b� �B1�h��=r�(�VF]k��fIPnl
ґ�%,"hk���X
v�f���J⵺ܱ�,�32����Y�
����
�l�J!G�o��{�	KY!�
�k|�u��L��7��h��`��=ڳ��=�c"�v�8�6f�h"T���p�6B�cW#�}~��|%}O�������tƾ���vjc���ܻ�Ww^�*��݇<%��H�F�i���q�m��|	���tTҵ=�*F�·f��d�f2S��g�a��d����w.�;���L��oP�z��ϼ<�ޱ���y�ܭe���u0���kn�&w�;�E�dΖ�Xx�S.�����QXڵ��"�n��b=�>'�{�Y�6!�y/�~�q'���@�hW'gI���&Ѧ��r��!b��8�p_�{|k�e����$*�u��"�3������˲-���5.�]b�RDb1���0ۆH���M������9X�V'd�'��֦�ϩ3��:L�ϻ�8υ�����a��UJf��P�j�V�.rq�X{il�2}��r.�LU��'l��cc�[2,�k�}�T�O��G�
y���2������M;��U�$�qa
�A����=
T����h�`o�r� 9�]��W;�E��I&,�D�b����|�)�Dj�d��n
�@JV��	2ňfXS�N��n��,.5��ê���cB-���k�=~��3_N֝��~���%�8�r&X�	2h��Æoyc+.�.8���b�q�Н�3�[���0[�Et]�q�ᓳ;��VW�&к��+3�Vхf1f��K�B����e��;�:`�$ɘ0�q����m�{��"NG�2&����R�/!�Ͻ�Q�M���xX�!k���^�>�����{�W�hR�QQ��
�����D4���������4�d_nW[��	vd�2fr�Y�}��k#A�{o��,��K}�=��὘،;��gIr��V�Xk�z�m̻f���jM�[����˞�t�
�-"�A�Ъ#K��W�@˔�^�_��i#X�F�B�`�O�� �H{e�vc	ڃ�d��ࣄ�����#��
&�jDq���9�<7X�7e��YB`0󚌅5N��ӧ��p�$�c�t'�!�����2or{���vҕZj������ː������"P�XBĢLAI�;&jE�&4��*�bـ�"��Պ�`��a.n�N�36G�\QM=���Ͼ4���9��Ǫ�gǈ�g�mxZC��ѿv�����hb�����/��:�i��r�8,��y�
�[�����2�	���.�5�<��7#�t��g���R3���N1d��xo��7hxn��8�V��� aG,���+8Ƚq��@rRA��fg.���S'f�Qީ^��ٚU����Է#U�+��B}����j����v���
z�PE0��S��1W:ƥ]��4\��@�TT�
�Ң����K���������)�L�Y`�����F����N�	�I��Fm�.�a�Â�sm�<A�';KYam�b]��2��1��)B��Z1���&�ԥ�l�i�Msa���(D�Zĥ�̱�n3�u�����<�������c5��1�B|A �|�}�YMU-
�-)G޻9���+�$�6�,���(�so��'�2�[�Y,
kEɡ��y4F���\Sh�
jG;C�,�3���t��m�Q��暈�7~@�/iv���8��遮,p����G(8�L9$PP�?��p����3#��5��~ϻף�>�P)��N�,I�y���,IK5ˤ鋻&E�n�"��^�]�������;{�D[�o3��"#fC�	�������_{*�3c���vœx{�C�G��S^6�9�۩>�����F4�}���צ��m���es	�,��i��Ͳ�&��V�0ìfvfM�	Li\Fn[]��`�Ż]�ؔk��Qa5�$6���2��ݑ�e6�f�iu�)�YM�`�U�Tj�Y��^sJ�p��X�����ƛQ�fG2��k3�C�鉂��pn�%�&,m���8�iiw��Ɂ�42W4m K��f#.��a?_k��Lc�����������[NGA���"(�v͙��غ��`���.I�.���b����3��q]XͰ ����* �-V߇����4��#���]Ȇ���ӳ�NN�]s�F�l��76V����-dxj���WO	(и}�{��w�꺫�nX�7�Ȥ�0{�{i��#6O����vk�%�$�.yI�l�=����Eݓ"�2���	�r����N��Z�*���d�}֯FJ4��U�#uV��U�Z��}ߵ��w��n�odȟuIm�6�����f�|a��>������>9���dr�.��#5(a�E��l�5����/d�U�)���l��4)RG"!�S��h��@��Ҩ�5J4w[��#=�nݟ�J��?@]8`	<נr##$��K�);?�v7ah��u��V\�^Ӹ��9e;ģ윞F��ĳ��7{\��kz������9o1�k��δ='dQZQ���EiDZ^}���U��m%<��vm^}6�4	�
3����\��4f�HG"�5�W�1����=^�~��7����-(]��$=���ר���Bfғv$-&2�Sl�%fsWn��Ur�t�;�F��6b"x@3��-�{T��_m�׭/�CM�d1�|�9�e�aA���Y �'	'fVx�4�C�«��cG�T4�K�b`*��ͩ�}=؛����1�}���y(
ez�s��lV��<5��i��GR����f��iQڷ5�U�W,]ܢ�t��&���Dx_�.���ֹ��gTN���*4(#PD����|��..�����	$�4T��N�^f�_6H�F8�����+����:�b׺VGU��g	9N� Y85ܰ|�Bj��� ��.�̝�{��t�6���Vo[^WeE���Sź(k�����v������J� ��Qm�5`�B"��(��ݚǐ	��c���%`�����,��f0�}H��fr��2%;����L�B��hܪ�n!w�̼���s�4U��~E5�)�����C{�����ֵ%��c"�S9OW�w���8���Eo#�n 0Ql#eͳX��>�[ӣ�o<?����B�@Y�,m+;@v���gm��`Z���y��nJys��
gK5��S���h>="���c�79���t�=�n�t��q�s���Y������&��8���׊S�W'<\���>9('��"���;��Ս�B��'R���6��jv�rə����3�KWwy����d ;�Y��T
n��T�X>��tQ�j�E�,�rggfd�X�b�����@7�Bφ=7��<���ep_�|�b�C���(Ɖ��Z�K���1��A��v!�-ӧ&m;pH^���tJk�`j�%h���7u��;���>�_������\wy�3�r̝�t�L ����;�B��3��tņR��-;�0��WUn�� �H�|[xV�)L�,���Yc��eY�ee��lZBj��Z� 2���sr.öգ����F؛I966����g�We_��ޅ����!����Ƣ.�6�C8N�Y�tC31L�c��+��rh�k	����ی�ЬU>�f�=-����M�ñ䠋g�~�v8�vk�-�Ol�"Ƒ�&���������#kޑ�@�L�$N|E�ֿwz��{s'�]��Pفǽ6N����P��9l�{4���`��0�Z}#e�o�����f�z�M6D=�����`��"�c�$�j�ӵ��b�u�\[�Ǔ>[����xv��WG��>�^꯽���[d����0�����3����m��j\{��΅���}"���x�}sQt�]���9ρ�#�>��:���DJ�g5�`񂔼�f��f�����]&Z�O�󏁹����a��19>
o��>�+#Cn��e�xL�L��Oa�^�r��X˯T�D�L�P[������?`�~1�E��ԆD�I I��IK���	�\��1��$�	i�$�I b��bI ?��`Ą$�� �PBHI!
 1$$$i�����!,`��H1��BI �$��@�1���UoU�6�=�+�t�� I m$	CLN�:`��hU��ů��dut �a�������BI I~H�����_ހ BJ� !$�4�(����"
 ���L_�W�4~�������?������IK�@���� ��G�'���4P����lg��A����3���?�~"�z0п6Z>�#����d����_����_���P��L~j���7��g����=���Cr�+��G����1��j�B�[+�P&^��⮟�l�&����!����e�A\4i5d	vnCz�V��馤�;�h��0o4�<����bz��Ю�Gٝ��p�C�rd�ۉ��V��%yg.�!�D˻ƒ�᝙Ե�&c{� ;��9tr/UrYA�ְW�s5otˇ/��\5�%A�x�̝!z{�0a��〕���΃��ɻ݌щ8�\=��wi:$��y��-�{�ynu9�2������q����*����Q!�m���҇n4��}�������&��SBΦU��s5��*'X;�T��q���W"2u֜�
����e�����B�'t�9�k����z��:����_vXt�խG��ٗ^Y�>�v��e�\{�W��@�Ιd`�+�����}��"���4q/+�g���vR�ͨ�=Ff�ø��{�'�{��Υ�q�Df���=���\d�N�V����n�$��uq��h3sc9�T������.��ސ��ѧ���1-%�Р�CdcY��a6}ƛ��fq|
�싆6��Kv��+洫Lz�1>�Hv@����@�tج��T2�ܪɱbʅ�pq����7�`n�GOQ�6�u7���+�gT��7yj�"�v��8�f+4h+�T͕Y��v�O1Vc�����<�C)��2�,ң���d��7h|��L��>S��9,'�l�1�.3x�y�>�K�4#ĺjC������A�X��͍pd=�m�Yx��t��s7T�zv��	��v�������nuə��GI=�~�uu���3h���s7sw����Q��-�]f��7�N���w!P�i�a.>8�eI�N�j�����ȝ��D����.R�[_e9û���ջ���MXÏrt�-���.a;�`�>5�6�8�GF���\AtPY�qmw_
gYg1<�#a	�;�5K3��1׈;�ܹ�]@�E<�h�x߱�:s=8wkh�!�Er�(b4�vr�q�Ax�X��1>Β��lڳsRxK[[ǃ�Ľ|]�1�8lRvcc,����(���pЏ=����다PŪ]#����p�B�O;�-�m��s07��G�I-�uY��n����s��#��z�\�=�M���:ȹ��L�aEk����;��غ�ò����X÷l���f&.�1�LA\�z+8�	T��{�B\o�^�ו�w:���`��3�oaɿ��Z(#*�W�|.?I-W3>q�<�V��4�����Mg{b�ˎ�{�w��ׯi8L�7�ǡ�ͅ�4��eKx-\�MQ�[3n�paΎNk[��:�j۽�:�Ϩ��G&�nc�]
�<���+j=��|th�s[��C�4��.niΔX&�v$�q��}�h��
�xV�쮍HT���q�'�~���Џq�T��Pox���rcx������FK��,:��#;��gj�n90���b�vw-�{��\�]��DH��ώ#܇�������;/T.�Fa"u�R%����{fc���0�����?t.q+�2t����*h�y7s4l<����y��O��/�A{���
�p�TDPZZJ�j�����*UAUZB��R��ii@ZZi�TJQE����DDDUAV��hQT����V���U�AJEUZEE
��R��E�)h)AE�ZF�@J�J���JD)�ZF��V����JiJ� h�@@JhF�h�i�CI h���C	CT�5H%-5@�U@4��T�E45@�R �-P#@"P��@4�
 �(5B 	M�QH%
SM)�!��C@��i��ZP(���Z*���j��*�h����(R�$�i	�!�I1	��I��hI��i�4 Q��J4$ؒm	4ēL��&0@�bh`�@�	0bI�@Ć�@�&�����@!�L@	4$��		�� �HC@��Mi��`&$4 Ć	��@� hC��1bI�hI��L@�&	!�&!�M!�CHC1�4��bLI4&!4�I0CM	�&i$КBiI& b@�I�&��Bi$�&�M$ēBbI&��&������`�LI4�I��hI�$�$�4$�I&0I6��0����I��M	4�I�	&	44�i��I6	0i%��H�LI6��M$�bI�I�i�I�I�	6	&4��Bi��Ƅ�C!1��1!�i	�1�M04��!1�Hi�M�MBc�HbbChI�$��i$�M	1�&4��$1���I&ēi$؄�hI���ēi$�i���ccI4�bC��@ؓM!1� �@؄�I �b6Bi �I&�&�I� l@�6���H �C`���cM�I�6�i 6�M�&$ i� 4�`� �I`	4$!�!!�$h!�b� ��@!�4��b1@�bBM� bChCHI6�&!	0B�LI�$�!!�MI� ��hB�&�mi$4 Đ�HM �`	0 @6&��	�-SUH��H*д��-R�B�4�I@�5BSUJ
i�!�� `��I�2�Z�Jj���i(i))i(��������AA�i��Pi�(��(��������J���� A�Q�E*�j����Z�C	���#�RIK�?�F���������Q���A�?���?����<�`��~���g�1-I$	/����A��{8��O̟����~_�?�����?3��>�t-W������G�?���~�I$�%��Y�4"�G�������x�����#���6� BK�RIK��?����???2�� \K��
A��������� I0iv�a`� ���A�G���ߙ����a�[��t��I$	&~0m~B���g�	$�$�����86�_�I�O�K�������?B_Џ���#�����G���Y�ƒH%�BBK��~���_�6���Bm�?�I ID�Ŀ��?��(������Rg�����?��A�G�.��:?Y�2͊%G����h�h�?J�:�~GI$	,"�oC��~h�f�0)�x�z����?I���A���`�y��h�	/���_�?�:�����l٤ _���P��(�&.�ɣ�������_��?���~`~���PVI��B��<�w����Ͽ��/������-EQ@*� P      T  (@       �EG�%�UQ@ �mU��@�      :�@                           �Ǥ|U��
H R�*�P���		(��*��   >� ����x ��   (( �"�F&���Z��;�%z�3������|����r[h�a�l���[r��{�U�yܸ}�v������Q姏;����� z��-�׫gW�u:=P)E$�7[*�meڻ�w�x]���� �ͽ���Ӯ�%�\�gסN��w�a���P4ޝ�v��nN��vƌ�Yy� ;���`���n�'���m�M��l��-���ԧZ qv�-��@��o  �    ��R �'|��!�] .Z�.��P�.X�֣�c�$z���Ё钎vu�4:��gZ����(��s��Qֵ���{c˶�Zۗ��tR�ݑ^@��$T�� w�:����o;5J�ֱGlֵ���ѥ�v�oG]h��Jty9<M����f�e�9��IA�v�Z�+Y\ƺ�k� u{4��(�%*Hw�      �`{=�Zҍ\Z��J<��OMإ�h���מ ��Ű
��m(���ݴ�����=����^ 2l���`v�Tvc�z
Q"��Z 
tQ��W�3\�J ���e�j��n�M=���R=4�y�I �9ݵ[$z��vf��.���������]�4��͕�kC'3T�t�$�R�_u�#�      ��V�m�}�H��@u�+�ԓѕ}{�v����f��٣���5E3zsӧ[e����Ct�֔=5םݠx d�R��;9
��N��BJB(( �*��=��x ɵ*�́֕K��2����+��@�� 6�k�l��jz7����Mov������
yQIAU*à     �� �.=(73^�݅�G���0(
�d���l�(R�P ��v��җ��^��6�*�� �Խe9�� ��`�T�$J"EJ��
����iz� 
l*� ���^a�F�taҦ�mB�� 2쪥Yj��t�jS�]�W-@S� ` �                          5<@)*��      T�LJUP      Lj���U(�	�  �0 D�*�R@� M�� %="	�U        �$��Ȟ��F��0i�~�Fj�u��������˃r�/���έ�m�$��PPW$K��~�@PW�?ń0SdE>
�����g�� ܿ��'����?�����v3������{{����:������0 (+���?�6�F†���������;������8;>�B�����/������O��>Z� �v~�Ӭt�~�u�|<�>��_������uv���P�}J�Pg7�O�����-ku�d�7�[��[�x�N�2L��עrv�F��A��-�6�pZD����ی�|;Ъ�-��1���n���B;�8�(����a��놦F���i{����AT�"*3w�4j1�m�M��ƮǺ��0Nךtx���)��~Tl୉n�������.���`��<+�����e�iҰc�c=:���O�>O\� �5�/�v��rt��x�L���dO"�ڮ�d?=c�.�y��==�%0��*f������~�����iB.�A|�ݟ�����"^}�߻�����R2�$duX�F
�(��/[xe�N3��>6j2���ݘ�ħJA8n�E�+���	f5|RB�{��wMvh�e��rf@r,ղ���"��znp��Co`�t�O�ݜ:v=���&���fgvW�p���kP)� R���62�2 M`����ʩ
�{$�CM�����w���:
b ,̆����Y6T�X.ec����Z6�:�9 F�Z.��;��n�ǡ�bv.�>{�n���`����/5v�S^�G�&�;��Gy˘�w�qX��ʔ΢JӃ%�6���4Q;��)��5"��ya�FH)�����͜�`��j��܀���`� ���Fu=�C0�;F-�@��~F�=�x��A���Nu9�g��P<���F�;;�{т�ˤ��uA���	�a,�-�d]�u�w�S��nvO�{��r���G�x����:�d!E������%4~!)Y*�^9���S�c�������e4���X�h/�g#�vL�����IC�l��)j����ݍv���W.��U���,ڮ�IA���x�8��0d��"��I�g�,�e\r7�[�]�j�Xᝆ��z� �z`g"�%��8^�R�C�I<;�o���Ҍ�v��J�zEF��,���`�5g>x��3:D� L��[[à�`j�X��{n�ǰ)�3��ܺ9��эN]Y-��'��`�rN�L/7�,zu��m��	t��=v��e�1�{�M�Z��*���[�|�o~�d��{~M!��hc��ɒS����k�S5l=L�˩Hr����1��@y�ؖ�[�rF���}��lǙ��}����~\Ժz�-�m�}�)s�PP�'o!�=�Kaְ��v��vf%��շ�}7�̧�u<�Y��כF'a���pc��Ė�עG�G�`��f#����l����[�R�H�n�����Ȣz0n��:Д@�޾���Ȩi`n������p����L�^�!9ۚ ���D��Ef�*�x2���3l��=Rn���8v�?�k �=����R	������4`â����J.`��ϣ�Q3c;ΜM{��s��2�0S�A$�c�q�ж�q��5r.YL�n��k���B.�ǜr 9���ȋЅ�^�c0#a�PԷ5UW�c6�].h<�Ǻ��X=�A�.ٔ���^ءKv�=Z`WD)q׻�v�(���c�%8���=V+NPB� 6�Ǉ��1�N}�ww:�ZV�Y�67k�U��m՞����s�-X}�%\�"&"�
���0~�#F��y��b¶u��؈��R�r�Z���]�9���s���-�:e�U��+p~i��髦�Vݼ�Lލ��bZ"l���lI�E�m����t�a(-�#�I�on��H��5+���}��򓳲kx�����j̹*ks��#�:�uf�m�ݼx-�v����ǥ�l�]��B�#¦ޣ���v�	��t�O���iG�R=��x5I)�ei�e��u=1L��D9�(�������Ѹ�e5�_ns�u���t��kmn�q��D;u�6v7�<�ln!&L�<ɏsN�vo���X��׬�g ��j�v�#��M��IC�y���;q����)�Ոa���x�N^mj�S�=]���x�[��&�oQs��N�������v�_r�p3p���B��6�5�l����a�ܼ��zS{����%��P���;Q#'b�xzҞo���+�+�;6s�$�EG�F*������v����nƬ�Q��Y`�	��>Fc���ZwWj�a�m��'=�2���z��T3�t���wE�]�"g�RX9�3V�k�&�lEE�J�#芌��w�PG�����&'�2)YT��x���L��F
�y�p=�t�7sbF��"'mKA���rR{Q��\��v�B����k��,���u
ŧ�e}��j-�{J�QNX��������s��K������P��b8�n.��$q^�茥������g��2l@E��m��nT�Y���	������#.������7D	�\thy��q�dYծ��z�f�X� )�Q��%h�Ovt܂�f醷�(�	k��OI�	ϻdF!��J�)�t]��Wm��z�v�,�����m��k%j�WY�=��;�q �Ј��v�j�Z��!e̷x�f�=�"x�:G�cǱ���sJ�yݷN��%'sV9���I%ת�vt���Fv�@�YBكB�����2��L�29nwN:7A��N�L����nG�cgx�yݳ��	O0E�ҿ8&�֐ۺ^/^4)Yڰ��c���W0�%^[�.�(�Ӳ�I4t0��n�\�=+��^��Xps��5�Nmfø�M�ݡI`@�L�A�>�6��G�����\�6v����K�����o.G&�b�wv0�5���i5Zw���#���%;)7����:En��s�o���'=�;V�Gʣz�q�}^sRɷvv	Y��K�]����.��q��[=16��5�J��Dݏ3�5�C��=`w��.�G+�?s�"S��4����Eef	Y�DV&�NQ*�S�U��X� ��4=��ú��3]�,��n�O:���r�*1=Ɓog3-�syn��E����ּ��ז	��eQ5gN�z�_Ö���qh�����Vُ�{�55�'�u,�wEQ�\����Ԓ-�	�/3���4hHLyOoq�(sX8X���9�;,/�Sz�y{$H%�7�v�q];;�C#�Jn#9AXgn1�5bC+�?����x�+�%nCܤ-R��vb��i�7��hO����el�f���p֚�����V<�<w��1��^�,�r-�\8{��{tbCp��8�u׭"47B1�L㓎��xVCf�#܊bo!jl3z&��<�d��M���Z�ő��i�al��ׇ ��j�¡�d�r�^���Us���6��f!%j�ڡ�wvK��<BiQlhknD3K[�A���Wpз��mu[ܢ���W��'o\O	~%��A�!��]r������͈�4B�'Uz���;KY0M��td?�3*�o��������ʎ\�0�ٷ ݸD<������];ŋa�k�ᩪ�&�]e�l�Iǚ�w�0E�os�>"�n�$�J0G]�ܧB�����6��y�V����F��S���vؗ���zu�B���z�GP�H�&d�7{R�ݮ��B$_��!v�AC���v�ubYvS�^wpV)�����yF�[�7�Jo�ϔ�8����,��3�^{�6{(˂��c5�DL�&�G�n���7Q:��k�+�<;9������]���zq��PMozEnԱ���?���wpu��z�8�Œ���p�	���u�/�_�/Zx��.�����_�Y;�]��`�ytl��]�wZ���6�toU8�u]cx�������zkx3�M٦�@������)�L�x��{����F�x��`���� �5����ԕ+��YѪ�q�+J���۩��GGX������������vD�M���k #w�,nT�RV�G���)�r�M�95~�*�wL�j��U�������Oe�ٖ�)��`|�B�&Ʊ<�ǣ��
k;Vu��f�t�d�67D���i�����W�	�F�:�hr���n	��*Ǻ cJ���v�Z��r��4f�����1.j�N�sQ�Pl���9���œw��h,��+gZwy�}ߝ�;`��ԩ�+g��r�z���kXNIN��זp
Q`��Zچ������i���PW��uF�n�Hf��O\���V>��&���:�X9d�v���ǥ�r,"j��Z�,��OZc:[nɷ@;R�^��9�4Ė�ٯSl|kԷ��}ѕ�k�P<-a	�ϙ��%
o2J�ZfGG#}8d�7Yqe={���2�2��]Z-�%
,�� ᵈ�C*�VK�k2��$!��&�.�~WD��]�Γdb�����y{;�not����;�f��fJ�oT�\{FG�,W�9�(��'ŗL)�x^�i��3a�N�T��f�"޴C�E���k*�j}�-2pəJ�a���"ӝ	�*�����x�-�˹��E����?�w廍�na`U,��.X>G
4d�J/-d[�H�(KZ 1@6j��y� /i�$�t��H�f�%�U+�&e,���]&�&�ˤJ3T���a��8jq\F($��$����m,��X9�l(�G@�w\�i-t�
KjF"�!��&ZX�)�Ia����԰}Ѥ�{����� dZi��o2�w8!�Ї殐#��3G8�0&������.�^.���l��g:�^����i��嵉�
,��-����IR�Ic�qɅ�����{L���!52�x:@���� Ca`���c@��0�3��1c���-�j�`�N��4�2���"FR�Z�U�h�4� ���dy���;q���8�W�nܷk76�#Oe���t��+�*C�Ct�dxł�cܜ���&h����ڶ���c1��N.��:1=�-������۲���6n,A�å����If�f%;��qιq�*��x�����R�R�2�Mݚ
|�3i3�B��Y7��d�u�r��ucPc���f�kh"- �X���APE�]�n
?!�v�G�Z�xA�up�< �f2�B�2�7t�̣ph�a��fau�2F��SY	]<��N��,��S'�5Kx�%᪄C�D�!1F�1L�b��Q	VS�v��V%yaVV A��!-�����x��
S�cfɷ��B�IP�"�@"JI���g�z��v軯[�w�o�x*^�ߦ�&�8�N%fLJ��jY�]�7�Dw]܃o�2fӰS�v��E3+1CM�I�,�Ukǎ���p���̈́ih�{���\��[�4�KtA�uCDZ��00F0������A�i���� g��	w#��$3R��/*nʒ���A�A0�87pQm��wr��탋�0�n\�4�+Z�z�5K�kmJ�;H����؅٩����sݗ;����V�� {ʠ.m�;������.8�7iܛ�t��
/)��F�k��;�7���yk<�}��qKPR�t0��**��t��%�M�qkcGm	�1n�'���k�q�4�<�$����޽ǵn]N�����^+V�x?���{���-:g:Ŏ\嫢N*q�Ջ��'N�JS6��`yG3��wInA5mˏkRlcpue=a��3���ׅ4�8N#Į���,�lw�~C
�������L��e쳬�u&�:��ck�E>��']�)�";'�8�\���$%�5Q�M��N��Ώ� up���
�8�'���76^Vj�5�]�%�����R3�&a��D-wGt��hz��4�V�
{�c�.���bPU+��-O4�'&���%�:�؟8v{�~x8d	�D1����NdR误iXa�:r(�g���u叉GA3`ʵJm%W4��~G;���$�{Ou��i/S�-�݉
�-[�#,��4f���wC+����cڷ jw56��Vʉ�JqY�X���"R�Z%�g3ymcj㷭m���m
���˭����?Ujc��!�&�p������b�뛊���\��M�5A�B��	LL���6�7�rf�5�8����M5�]�v�8�jY�8p�� ���`JY�G�陹E�TqE�r+�J!�$�C���-�c GX�n� �.�Bq�t���!���h���{����*���6��������j��HP����ȳLb��n;T��۬l7�A�j��L��+;vD��B}�xZ�O2V�`�TUZ6-��9�b��u/y��a�.�ym��@� $�iu^v�{c�����Uy1.n���=��,[�Z�R���$�?���Uv�����y��sa�ܺ6,�ÚФ�`�V*jBD<h���cH�!��_	ބ۬�Y�w.{�7�$ �]=�[��s�����#c���y\h��Q�����t��c������O�{V���=�����=v�x��Z������D����%����V��5n#xǽ�%����aW���f�֢Fq�Iy�)�Ԓ�lI�w6�]�an�Kt��7���ua5�S$�3B���B �1&Җ
��@���I+�m�7�߽�o���o�{�~?!����6�n"		�J��݄z.�'���&�����^��8{n��n����������8ٽ�/�ǥy��K�[�ϲwT�q���%3۶�˹�-F�74'�)�>:���{q��A�`Mw@�����w��<��ݜ����c�z�)�тq�5���x�dwM���s� :��vq���/c˺�2lJ�kp^���g��c�u =w<݉M�n�:݌u۱�\v�{rm�!{r��r6����_6܍ݵ���l�٫Mn�)f�]�v쎺�pv������ӽr�����X�q�vM��)�1�=�K�������q�,��;OLQ��*�{tWV�%�ҙ�y+��p�饀�&^��]��.M�[&ݥ���^9G6�n��8Ѵp��v!�$ݛ��G��탨�2�n��nnuEɊǮ����ڗu!����n��=�:�$����,ݷg��x��6�18g^x�0m�۳�sw=�C��P\W�^ܷ�\S��+��ݎ�,�u��͈W�8v^ݏ�6`�<6�\s�t��q]�8�mf�\q�׮�d�ӳ���-t��ϙ�ѓO��64v�I�ob�4tt��j�ý9��9�p�A8N�-��h�ιlv�;k��NL/F� L[��3���z�Fn���K��b�LGU϶;�R�l8�-�lj܏	��{lH�/Q���p��`n��arM�{.���0��C�[lu��l�.�;���v$u[Rζ^��;<�e�ٽ�[�Oz���C��Éi����n����3�r���c�w]��l�kv'�(���@��V���%�<dwh�N��7a�z<4�Y��ʋqt��;�0�sBܐ��Fx��M{nO3l/[p��*m�m��=[��-�n"�-�؎�i׶�S�):�A.y��G��V~We��<�㭝[F7s�/-�//^EU2�ɗ"�j�0q�
rƮ��k=  �)A�jn7��<r�#�n	��vɶZcpL$�['/JTf|��0N�Y����WR^N������y�z:�ν��Ϝ�����P�m��ݭ�r���8�I�Κ�=�ڴn� �y ��!�糌4�oI�i��+���U
6
^6�7�ٵ2�r�gZ�ƙY���0�KK��q���m��.��c�=e{1gI�m��s;�����v ��9ǁ���5n;F�-�R�dWg^���}Tz2�[8�`w9�;m��.��N��\7����kV��ɀ@zy֍w�O��ܦ�<ݞOnu����'KpEj�܆8���nc;6��c�x��\�;��C����۝���w9x9$������
 ��)�i���Iɽ��dq�[�#�힮���cb��F�u� ��^N��U�h������Ð�d7k�)���nw�.Mѭ��v{[u���g�����^�,�F1Uv��q痷[�Z�Oc�z��\�{���ӝ�����y|E�Y73����<��>��=�����V�n�'/j��q�L��w-��J��Ռ׍����q�=��N;(�7�5t3�s>p*v!��Z%e�u�����}�/hȹ�q�c�l�<A��\:.,�#��<�m�v�,��W�:9�i�1�#���e��q�'��ف�E�۞��ۣk4��,�W�1�nܻY�b�[��kg�ؕ�V��Ճ`�^?|�99��wFՌy�Oln�-���z�mGk��:m�cK�4Lq��q�2C�ϰL��и]��*n:����� �z�W:�qF�m/Fۆ����sU�s�՜�%��Y�wm�����Ϙ�]��#��G���nt��v.8t�1n��ܢ��gR���[9��Y8���q� �{8s�[�����;[*\�&�'Gk��^�1.�Q����k��w	���plr��۫�&h�b�L<n��x�y3�o;E�,묅r�>���pE�oi��k{b w�z�C����;���i�i'z7��A�<��q���E����ݣg��xn�a�Gnwc�73oƝ�c�z�z��[G<F۸;d�h��=1�<����=U�X�lx1�:`�s�mlM�<h�n|J>����=�=d���cy��O[F�=������'cVny���`�ο�٠�f]v��ٵ��a8ɺ9�[Y;a��yX�d���s׃s��.�\j��6������v6��ggF�;4x�{,x	�É�ѳ�l����/,1�n�n�k.x��/{�:*��p3Ɨ���Ž��a�θ���s��3�9�uE^�S��۷q���N�6��ۊ���tn�v�$�u����u�X�@�c�Ɓ8v��Z:���ɖ-1p�;:�ջ{l�[e!-��'v�~���݇��n�u�ܼ�������\[�Mآ�����ܻ;q�Y#ƹS�ln�JJ��)�����%��<O�����)�֮��瓠�x�r�1H�s���=�.�wN�[�{m�$�0a��qZ�smc#�c$s�q��'��K2�imr���L������&�m���C�='���6��q�p	�n�nz��lc��9-�S��(��x��{N&^�˩苲��~���;d���7j���vz C2g�\s��q�h�=q۳�rl쒰�Kԛ��ڦ;7����{v���Na��S����{uC웧Nsٹ���<����o�Y�Nz(l���|��v�%���s�v��COi9G�{������-<Xn,��ۓC���&�-8�u�����u�=�G.�'c�n9�n��-S�.d�`��c�=��څ��O��ݺ��.G	���xP�;E�7.v{+��2�[=���ct�G=�88ZSO1;��!�!cؖܪ��Pֽ)���z���5n��\���ny\�yN��J[��n��:��n����W+v1��|;t�M���F�b�!�
#�/FwX�J��n��y�;pd��#W)۞���l��Y� Wq�<n�\ە�v�<�Y��2�n�����2YC���Lw<�=����FN�;mۣ[G�z�2v�u�!��Oc!���ˌ���+�/Jp-k#�����҈*���T��W6������!;uqN���`��űq�@_/e����[rw�lU���(м//���l�V�)�W���l�m��v������z5�یo9 �Y����q�r[����.N�suŻN�M��mÞۗ�u���5-��yt�:v ��Sۓ�chڮ�t��������i���+̊gq���_v�^�f�ά��yt���0�ٲGs�},vI�����Zvk��7��g\v�h���v8Г�3ٹz�x��lFNzV�1�4���^���`\{<7q��[��f��������5�������O�c��q��cnx�z$��vu㇌-����kҦ��u
��m�ރQ�ъ�I�n��u�eո����ѯjm��틷e�)G!�a�.���n�k�jO�u��X,��n����u���:<��YN�4a�<��^L����aucq��\F _;�mk۱�����iOn]gx�;�Q�ݽ�n����-�8gd-�ۥ0S��j��'��tN���nة�n���;m�S�{\�[�k�h���\u�Y7nvMq�q����l0��ۜ�s�����7cv�:�M�k�t�66un�ۀ��v�z���;5�]`�&\Wn[;�u��ݴ��b%�<6�k�ke����Ȼ�.nNG�y�n�NGk�C>L�d)��2垃=U��w[��%rfˍI�&7X�yNݷ����۸+�ϵs�\�N��=�w>98|A������ݺ#<�/6���>GR�#n�9u�678�ޔ;]�y�P}�=��>^�kX�l�v�m!���.vͮ��63���]���l�[�������}�o��u:�y�5ڳ۠��㙺Ґ��s��SO�@{<ٺu����W\f��Xx�n�l���3��i�\�u$�]�LOm�	�w�ݻ���nޜ��5�5m�<��]&#
���!=p�M�;��1�u��N���Nq�iv�	m����a�ǈ^�z0�S���w	�M gY�n\���\��\�Y�-˛<�Fv&�gl�V9�qn��� D�r�����6��^س���0�E���3����s���:����[���8�.�v^#]�ڴT��\8�f�u e�lx�����uqM�/<�����[����"�W[��n��lg�3�����,ѹ�Iܾ�YK4S[s�1�����-n�v���>A�a(�;Ns��������}��q�V�9��;�zv݅x��g���m��%mh���[rH�qs�7c�M�G��޷\�:&ȩ%��.��Ů��읷����=]�c9�Eط/B=����û�;����_�&&i�#�8�nv�G�иخP㧶�(璫����k�,m�uŃ�1vљ��!��c\�g��r��|<�tn��;g��:��1�W\�8���I灱P΍ݲ��a����i{n�+�g�^P�.�7Of0�c���܍�^�����n�c�Q�6��[��m�d�.x�"��ۂ.�u�	�9��� ���k��[���X�o=�tѺ�Ϣ:h�s�YK��Ҹ�ֹ\�Y�힏{8��:m��pl�K9�'GP(t���ˇ��u�c��ݮGJ�j�;<�x�H{j��v'A��ۅz�:���X,]Z��zA�ݮr�wnvm�z��1hݻ�C��cg����<��u���Rb.N%�6;N�[�Ҧ���]���1��u�y��l���u��L���>7���6ێ9�v�gչ�e�;V�cm��B�����/Yr'�j�T}tW�h�w-m�!����Ft��l�̸	�/�[��!�|v��j��:�����)�C�n�;���9�v�;]����;!�<��`�M��ݸ�F�q�^DÎ���MMv�ü7j�������+nP�C��;�n��º.e�*��\�7n+���cP�n�mm��j�d���uI�m���f���ۛ��^�w����?PW������܀�j|����� �z�`�1���=��UA9�`�� rT_| �M���hhC�~hi����C�G$��C�r8�ܫ���6�@<�&f"<��S�\���p:�w�o�ޗ�6�Ud��̮�%�
t������n��K�,�v[T���9���X�����a�"���^��O�f+b3s/J8�<(��%g��E�]E����"bW��x5�>q	���/�85�s9a��^��*%�یh��E�c),��r�LzU�<A�	�4e�N�¶\HLͬ>qP�
O
�VI�q��4�=��z�ذ!�V4���	��۞�R�=��U���z�p-Ç�OwH�t�&j��9<��P��Ow���tB�wKGkdL��I���bA!H��._����"Jn�b�R��"�q�B�.+cD��`��Z�ǎ� �(k�����ovD:���`�ݝ�������n�d�Λ�;x��o16��|��y{�
���i�'Vǽ��,��K��01^P�w��Ρ�J��Y�.�p1��Xyθ;��� ˄9��=٢c�w�S���*@]��i�Zj��*[�Z-\JP��s�����+2�M�����q�|�9�;��p�f��W;�͗8,�@�[��z绺��Nzv.!U��+W�M�)��U%�&�EBS�F�Df�����_�-�>�����Ϟ�cҺ���;����w��=��Z���0Q�o�{Cz�~]>��z�o��]vaӆxjr����E4]�L�<��%�	�+�}W$��zb�$S�%�g�8�B��u�0�J���ya`�CB�y��1z�=ڨ�Ҹ�i�L�;SI�[�I*#S.R���
��	*ؤ�.�)����&6�]��.����ڳ�^A&z�,p�J�9��Ξaek����Z��{��pz�OF�$�瓼s�LL���c�罭�ŋj��Fk�ج`��[S����:j������G �S�7�N���i�u�3�[���U�rM��sž�]�yw��۰s.���W������¬��ٯv��N<0�z^�	�X�2�nFʶsIH�
�D�m���F����y�;��n���59V�G�8��]uY�b�g�p-�mEs+��	Am�:n��nP6�������Nc'#7k2�W	�2�ݯK9,��C���*�ua9�yS�G��1�T*�a�r����9��iN�����7[؝y���_k~�m��M��|��#�7uT�8�����/����^�Ǹ��1#��cY&x�{Fm���v5[�h�����9�ٰR&4M`ꁚ?N���Ιp��$?ov�g�5Ij��j�p4s�W=(RT̉���i�LD�����ֵ/_]��v��;Vw�oiJ��s|��o��#P�O����!�y����W��{rI�TDN���9'
�7=�#�=�����G���coh�{�S��� �˥�����*nuc7�w˞��G�ط��H*Q5{B���� ��2A�Z�d�wM�M>35��0{��`ɾ��7!����
���[��	��@��7��7`�F�_Sd��- ��P��{���j��!���]i#��U��\����u������;x�����nn?o����Q�%� ��mθ�������bsF�v�f�&ꯠ��ڹ��w����$k�6:g;"��a���"
伤�xn��-��$]AǑ;.��Fwm*ݡ�2���S;��gr3m#����0HVv�\>��_�|�)�Ղ^&����
o�Z�᛽��Fw��u��ž���KNS��3�ok4�6�͂=�[*�"��ebٻ�ƃw�'cYd
f��sI�&�l�7Ofɼƙ�V<	��)�F�b0j��3n4���N�	/~����=���<ԇ���t����^���rb��7{}�:������G5����O3'^�S�&!{o��{�v�
�qNی���:�X;��ʱm�M
b�OPH=�wR�k�yo��k�}�7Ex������μN�[������hrs=8�z�
��(|�] k^�h]�+w����<�O8*��:})�s�4����ڻ=��zf��j�۱ٴ�7�v ���p3{���_t����=!9�(����F�&�Z�b��|֒��)��ik�׫7�)�ު�+fP�Jy�L��)��ۣc�.��痥]v����K��xL��s=;�q�I��N��(��.��w�$��y�?rB����;��[�>���ە�v=��H��5j�9ot�ݐf�Ԍ��e-��I֕\?r��6����{�n�l ����,�a�T8�}}��Nͽ�ଓ"+D�8!F����;:�TԽўYs��n�V�w}1���E�<ڢ�E�ʻ}^��܀嫃����ye��n�����-z���~pN\$�_wq~�>���l�덌�J~�۷F(9��)��Z0�4M2w�-��e-'ڽw�}��
}�l��y+�0�uE�d����Qa�	Z�ֽ�!�N<}���-)�}/e����`�%�+��ߣ���۷��{�v��,�g�f��9ڝ7Cg��Kӵw�CF|RW��]�L}=X���p�N"��=_1�����T�qĖ��`��~��Ǘ���6����ӛD?�b�]�pzz���AA*N�A��zE�=��v�:��7My<�.�^�}{�Fw�bۛ�٦9�Ë��3	��U0�t�U�p���짝\mk☛�%�^��%�F"��lT�0T��fv�r�ÿ���?ӻ���ǚ�SY77�k�*���ç���wY���aU���vpr\�!�
Ou����]�F4�w�t{�����Q�`�s'V�*u�/vtN�wj�UX�d��pۊ���Z&�r�e��Q����2�|7����1\>�ꈇ��B7����\�9�����#���,����9��ey%$�:�,3bq��;��xu�4C\f�/f�Xل6�M'1�Isȗ��6�t����{���<�G�l����9��o��4V�M�鬌U�M�0����6�u25_yѻ��ݶM>��mP}��6t��w-��8���36���y����.��٧<����r�o`O��ҥ}�\�ٞ�5�ç�s�t3�Xo�ݾ��0i��g��I-Y���{e�d���á�f��2N`/x�&�wX�?��po���iL�3��h1���h�!���=0�J�X��y�
�5���w��T���2�.[��+9�?]�Go�K#
�����<��0n.�VS�z-G��a���n�i7�]�jrf1�4����W�N
��A��v��}I�H,o�Q�4`ח_�eV����R1�)�^ӌ���f�<x�^�F�K�A%SH=y7����ˑs�J�N�=��䳚�A�^]*́������ʝ��Y���1^��3��-��
�;�������w=���me��P�=^���H������D�q��7�`cX.���^�*�9=�D����Z'���m�hW��Vn�����%	�$�[-=!��cTY�kXʷ�4�1�o�ء���c�B3�����S���Ujqdl��Ӽ3�}I�7��	B���4 ̪;cD40T�EjѮ/$����}e�j��I�}�a��羽ݞ��
��v�>Ùc�(f����X�7�/�w�O=���叺���@W߈�|i9�i+�cwz�_����{��{�yw�q�๽LM^��|�w���۰�?2�(+?�'�o�zzy��̼��m���ȧ�n�e@g ����8Q����s�x{��ms���k�����(�<���l�r��m�����'{�E�9��vxa���k�V����͸��v\K�,q�$���ӗ4�{c�[C�p8��mr+m���f�1[��t;���F�xϛ=J���yi�D}���t�8��t=b|&�$��S�Ĝ����s��&C{kwn�y���;x�mۮƤ"�95���wEcv۳��KU����5�x�M���G.�-�6Æ.�l��gH�^���4VZ:�Z��Z;cs�/m�st�K��]��ɖ�
`�Y�Ax��3˝�7c}q"�=�7f��{f:7rf�;��f*�n�5����c��6��D�Fz1\.�3a۱�n����&�g�ck�Y�۳quD]'oOV�.��t����x�nw��dNt8�*�O=K�: ����Z��V� ����VF�bu婁kB�N�
En���n��g��8��U�	yc'+�w�[�s�6�n�B�;��ە��=�;��C!j݁;�=��ں��ۜ\�y��c��d���ڱD�z��$��]��n�_y����5�uˍwH�H-"����=1�9����66�8��Ɯ���X�:yۇV�����¦��ض��mwc�'����u�3l,���뫶��jJ��յu)��+n�޷��WY:<�v��۶6�-\OWs=�l��dU��=�"�n�����<��lSډŞ���3���Y�GAד�r�E�b��x�<hy(u�w�ⵦ9Nđ`z�9�˵�9��$�4v�Q=e5�i殰�]nXD�+%�ȑ"H���\�^�6�x��3�G��F�a���lݸ��1�P@�5s�&^�n�x�pv�&�%�]�x�=t�7�&���;����a�]��+&�k�]Pv���7����ۣtp�v<M�cۊ�\�ݺuv�\l��^���t�p<�:�]��{<u-G��qٹ�[q��K�[	�����
Z�@�8�eA�U^e]q�K��Dz�m"R�;C�.����w�"�(u!��{��iO;�]�]Ƨ�k�!�C�)�8�ԟ����2v��T\Ԛ�7�Qw��_j����{�wn��f���MIn�O�u��h�F�a�C���q�i�%>�k�n�L����"���[����0������jY�T��뻞k���D�f�#�h͎�0����۝�ݔvn@�����ц�Z�Z �c7o3���Cgj�|6�KsѼ�ٸ��4��}U��ié�=����TP��/v�׹����U�s���z^���֏��n;?.��m����;�k�0������qQ��ŵ�����"�.��0��O�pKx��Q�'�8�8�c��s��쓸��cu[Sk��>N�-��!�t�g���FrZ�	��z���Nh�vKum��c<V��ٙ�M.���^\�G\t(��n=�ۨۛ�8M-�<a�����R��v���ɺy+!�ŝ��zn!�z�$+�CV�&�bNh�c!�=Z�C�9ܩ�Y���������˦�n�d�ίҽ�­/yQ�.U�7�k�QU�Ϥ���]���h�L��ܻ�NNɷs�S�<oc�M�Tx^�+����� P�@�Q�1.��3���(� ����U(��*tJ��:dט
s���޻���z�

�**��ФEDQ%EUU%Q	J�QAIM	TR4R5@[�DIHDP�R!R�-D��II@Q@��TRE!BRE@��4�P�R�45M-%(D%!HR�(�J� P4Х4�Jд4��M$@�1�����ih
�(�%rP(J�bP�Z�
Ji
j��j��J�T�R�)
�i
B�B�)Nw�SBRPBDRR�	T�Ạ��B�R� SHTR4�AIAHR��4� d+u�d+BP)M	M �R��TP�M-*�P�4R�4�-#HD!JP	E$UJ%)E	@�KM4�4�0gR�QICB-R��$CM"P�T��4RБU%�KPT@P�-!5T�R�AE4��P��-QM)5�&�q�v\̸�F�[T�Z���((�)*�i�(
j�����((<,�����"��(�H�"(��JF�*��Z��(��`���*I�����E�B
�!D����&"���& *������jj]��DP�SG����P�R�Q�PR�4�m޹�7�8�
j������"J���
(�"�b�� ������(�b����"������\kSE45CO;�-%1M4��dCKQ51D�`�EoeMPD�T�BSEU5UTD�Xc�E5EUE�U��$�)jb��f)�����(J	�!�ف�]�EUT��Q����QQIIy�kS4�I�%15�--("����������&���T�TQAT�;�EDT�UD�L�"5���r\��!�cs�ƅiR�����v�6��(k�(���¦������|��$�ۇ2vڢ"j""���	�a*��uс����h	��!띳2t&�Rs�����JH�Ҧ�jy:�z=�B*j "h�¥���ѽ�A�)�P�1s	ݨ��2$)�*6���3V��&��
"(�񲈊�#|p"�*����N�9\CKKF�����.�䘗��Z��*|BSN$JUh��;�{����OQPiZ*ܰ���SSP�ڲ�)"b�j�˼1�" �"
^:n��X��y�N��Ֆ��)�DAޖ��"�bF���f(��HF�Ut5�D��L����l2��j��i��HNjM%��2QEL��51
����-�uyXZ���U��.s&��h1� �Z�h�ٍܘ�"Ҩ���A�)Gܗ�u����0�)i'�dj�i(8��i���F��Vf@�w�ɕ�=�iZV����E)�G��R9)�Z�J���~�����c)��F"��}������]������[��]U��s��� �
��M�^Fѫ^���:b��ӹ+��/���Y(U���H����]����P�h�lbDH����;4M4o��dm�Z
5PD�O��5F������̐Z�����i�i����"ѭ������WC2���鯆�!��/2+�������w�� һ%��e�%�F��U��qA1IK�ark.Qi����R�b�6y�l*&�8�Ȫs@M�;���|���`w�g+ٯ.r�AkI�M+�Ȟ�PȪ��b�[g<��EVZd��'P�:�m�����Z�Ub�<ƪ��3�m4��- P�p�0$Bă��S��Z<��ѯ;לk6�rDo R�/r�R�U)�4�Q>;��x��Z�/"ͦ�y�i����)C�$�C$u�u�`J'������A�i�&Q����P@��"P-�PT~+.���u�n�g�0ha#E*�r�� j�����J��Jy��ThNz�mm#�	�J� ��nH!�Sǘ�k+ō���ϧ%՟���v@76-�EH�H�Hm'2���_M����|�*�m6J����$�D�^ �� ����;��C�'%B���R��C��Jy!6�L�u;ks�t&��#��6�A.1r�6��~v����7�3f�tUi(ZZZ��!��(�Ȇ@�����@d����)��������k|�3Z�+&F�H9/;b�����Sg1l����2R�C�����8��v��-�SR%-t�NІ�'>8��b$�#]�	�8��u�\�)2�
 ݔ�%@�U(�ω���w���nF?as�;9�qkry�]n����	�frb.p7X����
�:�c�kf��5Kj�UR����CH��i���Jj��)���Ny�zDj�IT��o���@64P�&�* 4�e�-+5���k����K��&�]��F�Rh�2���v3	�و�P&B�d-'�;u��s!%�p��YUUm+CTu��Mc�mW�*�l���>�p$��
%ᚐ纱w�}�G��6��8�z�N1hD��d��ϻ\��S�([�n�o�Tm�����|H�=�/1i�������4ij��X�]X;NE�!��Ay�}V)���|"-&�]E�ˬ5P�C�E�^�D0^�B���E:�ؘ�<)nN���3:3w��s���;�id:����u�ED�������׎��7�]Z �	�g:�Yt(������*�k��0
"���/�X��Qd*?RZ���1Z��fT����)5��ݠ�b28�(��6��<���-}q�Ʃk9��ݪ��&�>j,�[�������2�)�D��g^kD }�~ �Ș��=����Jb�eI5ʇ0���+m�hJ5��w5�dȗ���n��W�t|Х����i�hk�cCI���,w�ٿ}���%��%O��"���x{+�&ו4��)K�R���<�.LЩ
5&z/���5���)�"e�pر&���rFl[n%j:nW���y�{h�hd����/�$bt>j��j�ƫ���YXҬ@�4i��E����ᯯ�W���xcFn�{��Ô�|��m�\"w���NN�"bLMf6
�j��Gh�0����k�K@D5�6]b�Y�{}���G�.�O��k]�ѱ�%"Mv�^�i ��c_	X��Qz��7칼>{��}�JƲks����3ċ��z%m��A�k�tVڭn@���H��G�A2�j��FR�x�A|�=���:��	\��FJ�T"��F��ߡPGb���+��Ŷ���\_-̓q
&�ft3]�>�	${|`ռM4����{�Ɣ��)����H7�h�2,U��������<�w���9��s|�E�
�{a��(�6#(Gw#}�#��)֓��,��V};���p�����yvqGآsVL8��q�(�����`Èa�Pih�i��|>�L�67�-GE������%����0aj4i4��z��U��b��B���c+�5�/f��v�ύ�A��y�z`��yO0���\���Q�QS%��6��ƺ\	�n�Y6-O@�/=�m�r��Y�PX��HcK����$S�WM�C�HV!�v��
���B�m)5��Os����c<�`�` �*�$i�"0b����Abh���0L]��^j4b�pk��rk�<M`^�/MD�N�cW�����ɴ���B��" ����{-P�{ں����\x��*�|�qO���Z�v�,�2+_ZZ�ս�X?�Uv����@l����J������t��<.��h���|}�.]���"� o�Ϲ�'��I�chtg'͢�k7!k>Dh�?VMۿ9�z�F5g�оt;�$ yZ���H?>�=�✝ܷ��7GO�L�c��-��[�+E�yı�~�~��Z�_�щ��[�>/N��4u�Ī���"$�Ws}$-T�凹�A�Fa�R�K��M*cL'J�|�w��3}[8Fc��n���C�&��s�s�`R����g1L�hb��a�n��m�u����mgV�L=��kWS��Fs��n[lgg��m�.S8���X+e �;	�ם��w3�lU��pvc����S��	q�f��O;k=�v2���OXӑqMt�-�9h�lt�D�	M��kb�nֽ[v���θ��؝tݪ�T�鳟C��ǴEN���o/J��K{klV�Q)	��cR��z�j�-�Q{g<�!]P�t��^���B��'k���ru��n��;[r}s����m!�f��k��+xV0n�*���7�^�f����\~���ykO$�����X}ͽ�u��ARh{��j0�{v��\�6w��ۻ�����Z��6:�X��R̮}N�����>yO�A5�A���Mr��ݵߓ-kG�_^���� ��9�,��1�h��>f�
EP��G�-,���r*��N,�ib<E���ӚG�����x�1��3ej ���'B��`I/8 �<��g�2�$�K��7q�^ߚU�=X��v��_�\���`�¢C�d����X*�e���O_z,�'Nv�z�~C�jض��$E �!_r����HABK�����tO�V��q���<}X)��h3�{�s�I'�=�P"*�RC�A�ސ�����{��a�����\\*�R�vW\vօ*JW�j���;F���][hxN�O6�����mM��EU���8���x�ۇ,�\_�o�I'e{��@X�����GrZ��^!����
�bh1� ��NЅCE�!$!B�G�|tZ�8����nw;#�k��#>����nN��f:ۯ�QW�t��}�vv�b�����xY ��WS�)�P�䁒�r�H�� �"���Ю�g3���O>���!
�!fk:��w]s�*��1b�s�Q/d���Ͼ7�(�:"�K�Qz����fV���Z�<�2�6<��\־��L�I�jN�э�V�2�]g�x�\~�Q�.���s�V������g��˛��UvHS{I�K\x&���֯��i��^{��1���C�1>�I��w3T�bnŰ�z���ܤm2������}ՀJ�{�N�jP�@��+Ĝ e�	Y<�Y	e��X�}NrI3��:ӺN"��%�}�y����a�+o�&�|�17z���=�#���/�-ZA;�zanE�^��6S:�)\W+�-)�{NY�!���k�<���F��GmrC$,*�$�>b�~,Ǆ�]�;��S��mC��5v�Y[}���P�+����/n�ӽ�����˼�+��SMq;R�}���'N-���4���`����������% �8	'y�9����N+HQW��P��\'D��_���Ϙ���}S�@ŏm���^���d���*-�a�=�u�/gu@Jg�|���G���p���~4�u�8�h(�*� #�W���Ԡy ���D�no>�1��ޒ<��)�}��I����5U�
'}�o����W����y������;N�~���7�Oݔ��C�5t��sT��T�e�nCSO>��\UGe�E$Ms\�ѡ��ύ��I�ֵPW�_�v׽���`}M}a���m���>��D[���_gJZ ��cmmN�m-'�'YbD�5�#j�5�ص8�����&:/ϵw.J��6�ɱ]��ԭ��o;ܝ�s[��&�t��r��S�:!��q� N	41J�Хm��*ǳ���9ۜGF������5�P��"��*��؟~O���8ӯ}�ɡ�.��j\�# sw6��	�2��Fjrqq�^,�S��� �J;����jL����5�ժ-�ڹk��:s.pm�E�� ��<�(fy�P����2�+g��M����_�K]�i���!L[�~������Y�����Jbrߜ@ �/xD��j$�jIK��$��B��=<Q�,�����K#�]�/����o}Xψx���,J�b��T� �M������C��Ss{�s�����%�V�;Q��21��s�aj��KSB:�-	=,��1���b���{�{��kږQ���7�����t$�`#�����ũv0O��8��4�|�.%B�M�O����X�D挫V��̬�����0Bq`2G5^\���ND�IG�,�yO�ĕ!	$������;}�x�e���\���SnvF�<��2$�wn��t���N竟�vk�l�&�/3.0�r��k޶*H�4:�3�I�;�2N	�K��f���WJ��?!M;u��)?m:6@n�����٬��g�g+�u��
5ϟ��[�ͻ�V�xn̤�eK���׹�^x�9~�.8���o��,�eb��n:�:Y�%�ܑ��;%%y/�S.��ɇ	��j�hf�RIv���U^3V%�s_|sCwjc���c�O����~w��J�=�8s>�ʸ��e3q"i�^����
˺:����2�H�>�W9�gp�	%#U4��k��sZrI��ġ��G��Yur�J�XjD0�4Ӹ-�x�Ԓ��p�oﯚ�4�gD��]��N2��ڞ����×�WP�+fe'vE�%%��u=w�.\�R�&rBg�������~:8�������;qr��]I�m�uof˝ۘ=��޺_��u�3���iLl�l-l�Κ�OԷC�q��=Fp��b�Mrq�	�W��u<���N�lK��nݻ&{D9�o�_mc��籅g�݌q[]Tih'��r3��n5�iwm#�7!]�#"�����sٱ�������㛭m�i���?wޗ펳�r�Ωʧr	n���^�(�s�"��>��Z�Ό���h^W|:8rc�3ц��WS����O+��ld��V��Ց�M֮��l��L\ȌS���m���_��+zi���E<+R�_Y�l[�*���X�]R(�����,Zw��l��B�>�n�H'e)�`�]:�v�bFO��H@DFz������à��;�fT8�K������v"��P�5��> �_���Uh������u\vܙ�������8���Ol��$�J%��4�p�;!q;QcO�ѵ�Wy���˺�8<��� �	$=�O\���o�L�������w�$��7A���������X��c���k��+VuY�-ԛ�t������iG��;Ň���@�^��fC��?Uu������۫O�:�ۣTj���Z\X]M���p<8��v�Hr�n����/�C|��ۤv�Q�?*�!��_�_+�˓KJ�3ޅ�����D�O�@sǱBǰ���u�ȔEi���~�z��b0\Cl�4��Z��݆AG�/��Z���Q��l.��D��|��T��+wX��[̨�
̽󍕷m���CFr77u ��X��ۿ��5pJ��c�*J�#�`��GO]�>KO�xXY��������Q5TM5��5�>/��݌�Yc�HC��{��͇E	�'�{�&��12獃������ao'���oU늞��jCR:Q�+@� �θ��=�z�GO���Q��X�;��D�y�znb���2l�[8{��._!^�pq�VDP��w�7ѧ��j���,��͊b����G)�S`��R�\r$L�Ns6I'k����㰮��ɴWE������-�	�U�,GD�d�IX�������D�8���畆}|�5�+�5S�Olfg��"�S���7�� �޵]aC۹w&L/e�L5 ���#���s���\d�~P��t
�y�aq��uz��{ʺA��4��2B�����#x/���k;���p.R�s �Gz�fD��y�/��r����?V�����edQ̎�O��x 艥�*��l�K��Z����\���f����݉BF����:X�=Q����y�ھ���D`���䁚�bσ�h�lg���Ur�����QZkSs3e�J�!	��1�����@������Ὕf�4o
�E��Dݼ>j���ǵ
ܵ�-;��bw"�5+9��1\�b��Jbz-�k��%H���7^��p��k^Mtq���ؘ]���=��`�5��ܥe;��[��\�a��v��S�����{�"�VsĆ[j��<��Ov�n�h����ݻ���Q��O��ݦܡ`W��~ޫ�͘3�{��~[�>Bv�	7ۂ\t�bjΕ��wR�wZ����#V*U���v_n��ڸ��zv��=ؽ�'�)?1�VЊ��쬒���4�6�'I�
%
3!{��3�Ў�)���sѹ�&*t���X�_#���6�[�5���8$����%�{Td��x������L+��FTȺ1&b�3Χ\3�qcB�=��j�o��v�ɚ�]*�`X4l��.ڃ%����z}�
O�V�����/���Ƣ�ت�q5�.�l��P{;*j���i�8��ZI�q��GL�OD�q��YV{�3U���Gx��o�'{�y'j1f��oxM���7�$���;@��Rؖ���J�k���d#݁�*���b+�t츜��X|���R�&������3wXȡ��Fv	{���quL�2����D%T�/q�ґE��+J���G��`���ڽ�.��U��#M�u[������&��kȬXh l7�\F]�/sc$:�mi��Έe�:Ą��b�
�����7����q�G���ض}���lڜ�o;6�B�KK[wp֐��6;u��8���b�30"c��e�%��;ү>}�>��>jrX_����8+d�*�V��<�Rbo�@�#:�*j��j�8�J�s��d�*��;���t�*��"�gr$اӕ�]͖�sz&��Oe�N\1�_5@�"oueT��+��Ŏ��SY]��7��3MK�M�ͩIm��\�<_@��Ն#NI`�{�0h��u��k8�ljl �����ϧ]jm�{��_��3���ze����U��]!j��1&�,�͑�4!e׼4�G����,}�� n��!/E��K�|�my��+*�cy[�ޅ�L���ޫ��ܧ�xK�fj��Mf���S��X!�\�So�I�G�MG�O�"��{!��_w}^�}]W+�ca������u�F��z�ߧ-�1ֳK�Midd�I։�o+fu�oԐ!�5Y 8!�����+��h5�P��0߭=�����5�l�$���~��&0+��|�B^M�}x�7��s�:�C�&��
�m��!&�*�f��d"�ԉ��A��KJ�{t�X�X֎r������eA��Sd�(Ϭ�^�$h���;6D�n4"���|���S��,�S���\ԗ]�v4�[�TzskG~ןQh6�����cڹ�u����}��L7���yz��l��7�|{�x��*���!����\qc�~m�p���e��Z��A" asn���I��}�޿B��[Z�{�n����r⮎S🟲�)���Y�Oݭ`4��u]�QX��H �o	<�(�����#Y*.Ɛ��*��ʵ;ũc�`�¥D�]6?�<�Gg���_�K-�̩�h�t�@�k������|����\>YP���z�Ϫq��q������U�5�ħ����V_��C5J��R��������]����ή�s[�]��`p�����i.4_C���n��o@�軩}V�N���=�c��|��p�N�劮��E�I�p��;r@��I��y�^}�j�c^�F�B�{�r٪F�JZ[��\�T!��v��C^޴���p��Ѻ+��9:�V�4M��@�nHE�8GSra�h��h�J��="<,|)
�C�*�����۲�|�0�c�Ma��%�uFm�κM�C����y�6cc�7j�5;Ƕ��.��5e��p̵5H~m�U�*Ρ�GE�jYz�a��71�#%\ԫ5>9��Q�����h�Wk��v�k��!)	�j���pk�!��3�U�ϓ�ݪ�+n�h1�������>f�,�&|}aA��k먌������AR�ʺ��ԆԳ��'�?���h�;r�x5�JO�ȟG�aS���/9x�0
kH"�ϻ	ߗ�b]�X�ʥ���YHrF���͜���^-�s��y�B4������}��}�MO��,'���dd��Ndve�-a�����V���,M���~����)������|3�9�fH��SU��`|W}V��3	��3G��������	��!��4��*8�I}�Nu]�0�K����`j��Zu=�®���e)��h�{p˜�{��+��.��a���[� �Jb\e[E�g�,�Z���m�e#��s�x�^V��\M����W)&T-i`aO��RF�4~�����T����Zk����	Uۨz�tH�F�^��J�U���U�H&j��a�j���X�b;G�1���yms3�Y2��⯃nk�~ჷ �"t����+����H9��j�xDVZ���j9=X�,�7y�
��dDޭ����3M�P�0�.6�U�=s���Wd��kXkSq��F�N�lbwVT,���������]ڷ���[f�W�{l���p'C�4��v�\�LV�l�\닃�=�mmـ�95k���.K�!����WB�H�v��۰u.�Ս�rRx ��g˯v�cz�;��h@�>.{�{\������U�n6���@�r�v��X�׹�@edQTұ��������~5H��\�O"���T�nXّ��ҽ�o����Q�ݲ�i�5���]�,\�%�ѓ�h27���	)Y2�P��}5������ʢi���G��Xj��6p�0�~^0��C�)�l0ެ�I�},�;�a��ӷ`ٓx��0`ԙ��.<^�q�\u��3��΍h9�w���xt�I*Pq�S[��R}��~��K�\��JF�&k�?k.T��Ry�gDԸǢ�v�Q4u����'��0}��,�gն��sLU�����,sN^%5渁��z�����I
�}�U�
��fWxaG 8/!UR�Z�@{���=$�����$�%r���CbD�����j�++d+E�x�=��2���Y�-,��w~�u�Nf���e?IA��u����i�)���2���0wӍi��4�f4�F������ϭ�j�K\R��ʜɋ�%q4~��������R�}�w�v5��m�Di�'h;�tV���b�'1�r-�u��X$ـ��}jnzz����#֫ɔ�@��SMU�~׵�=,�2Ʌ�s9U���;Ι=�����0�os�`�n�`�D��>�|j�}�d=���~jW�	���F�5it�m+�YI�M�Y�W�����܀�2@�R}�ǻ�q��i"�79mn�.��W:��t�ə�U��^�t@�u�tF�0����~x�̮�BO}޶��Ĩ�{�Vi:ѿך���-2� �t��N������CCėX؉�e"�߈w~����m��J���JV�%?�]�Ut|�j���j*)�v����ӈ���ڠ��{��y}�$�)Z?��+J�5�uX�����r��m�nLu�C�2�Eͼ�Qv>o���������f�G�qq��y���Y܏���0Tx�pL��r�Mvm�+���q��D#b�!���-�����Ts&�4�;�[��G� �1Pi=uLw0>t���)��cKV�����++�,��|���a�ҋ}N���6F`��'y��I�U��l�M<js��o�Ĭ���Ϗ�f]ܤYTd��<��)�b�~N��~����&ڶƔ{S�>Շ���Z?j���]6f�W��C�y��߽f&�����=B�}�ֶƌ�85ߕ�����X�*ԇ)-��&��R㲠$z�m<ז����>oS�:�͞�������24]n@G���ZQA7�FCh�U�D�BC����@$��:]_c��4�~��rΉ�Ѳ4ck���Ӟ<�������j*2�[�)��WQ!)����_T��u��I���M!���9�zg?�Y��:��j���.�IfcǋۈcEmxB�fV�{^��a�;6\4%o�8_�Y+T�wP]�3�Y�v�E���Iϣ�D �Bz]+�][QX���+��۱=u������2������ ��N'�:��/�^6:W��)��Z�N�J;CΩᒖ�,��]!3.�j�������l�'�id0��<n_�}Y���J��ֺ��gX��i����+�}͇��"�*�|RcmN{���u�C "��7��~`��%Ҵ�P���+h��Y�j��n��u����ZA�s�auG�Օu��q�"��P;����0�ac�V���i��t�j��{:�h��#si��[`�6 o��;���!����f�i�&=�oKI�fa�PP�5ˤ���k�t�e>������F�P����!zw��w)4R�����4�؈r����� �S�ڑ�p�輠�s�Ո͘l�f����D�γ֔-�L��.�pv�Ϧ]��|yh�L�_<���y�D���'b����s,@��-.��m�敚���lˎ����Ǝ��l7Yz�+Z����ι�M�e��x ��#�=Ӥ"���vi��'�s����hpweƬ'T%�(!Md	z��k���s������Z��y�g\]Ҵ��%2���{_����Ԏ�W�z�+�9���լ��ˮa�ߜ��q���ݣ�8n-e��NB4������@���~b�
����'**Gt��9�[1�4wa���]J�$���nU�5�J�a+Y-7�q�h�a%#��eϮ-�S]Vڢ��x�M�����O�;s-�ѫ��[hRB"Ym�H�T265>��?��O�@�N��B6�[ks7��'�(���_/T?$��W��>l�M�:Z��F�z�	�i[$����ev����s����N�#V<��'��o�ؒ�m��j�*����^���^0���p��g�.��MI��]](s2���~�Od>�\��e-�<�����5��"R~�kK[͡a�5u�� �b������eJT����}|�=��x�i7I�LD4�o}�-˼��rd�����TNT%*�)��/�5t!nۤ��$�t����	�%����a÷�GV��Q�P�c�-wkb~�fB��l�!��}겱��l�Me�U�����Qr���ˎ*�I��A$�}rc�}�3>�z'�_)������ n�!)e�2��D�ʷIU!*�.5>!v�]ߘ%	�}�\"/�{6o�s;/o�m��buA鮱s����WS���c*º�5�M�̡��2�MkI�;vb9�N
�?_|� j��K��1QY��eYr8>�[�l���r?��3md;�=��ku��.����9����K$(܍�[Ǔ�v7q:����qE�֭]A�z�3H_?�������;�jZ�AԜ�?v�,oOi�&���D����G} !�x?�bא�VIf�P�'�{��\$y�l����9��]{f���]��)6v;i������o��e�5;�j����~�;tR�j�L���5P��Ԧ�B��+wQ5%.�d������5iVP�o�d+ ?t[y{K�NS����GB@�s��R�.)��kI�d��JMX܍f��n��po����M{9��b)����]M��{�`/�W͂��S�����d9�ڻ��'���1V�(���6�F��������WjDhY���o���Iq�z�F�����&5?p�+$?W�iȪD��l2JY!�R~˲��$�_����ߎ|Rv�_lt�5�#Z��#D�:aۯ�U}�ڠ�u HI[`N^�l��Q��p���D�@�t�C�����x�)���$��E5����C�ˬ����54�NSm��mY[H/���Ȕz#�A�o��CK�Yj7ہ� .#ٍT��.�u��}��&dKBF��B{^^�Q"��R�˯`��=��0
ar`����e���ܲ�T����m1�v���D/���?f�cJh�ѯ�;N���^	X�BkFe[��
o����W��[O��`���耉�-�ǎ�N�S���+�_����ܱu���F�G/��8$�/���0z�w?ss��d�q�Y20CTj�
�;l���/�o�'�kWhݫ��6D� ��d����'��7a1�Vۈ��:���ø-X�莽! �л���b�5��%�]��6��r�d�sg]��֌�h�F$�[���ID}=�7|���s��l��WL8�;��q�6���x�v��B�㰡�X��������0U�${q�$ԏB��n��qt�{'DB~@�����>�𲎍�P5p���KWy6��ɭ���~�l����}�.�΋�m\���Ga�8�-�e���:M�2Wqw��zL�J�KB��5�{�)���!mI�oT�����W�3_�h,#D8ok%Xf����"���[P��'��fe�<��������ԐgΞ8GȄ��2�bAl6ϻ�����I��cz^Ϧ	���YZ ��O�أhe[ ���a�=�n����{u^�	'*r�Âp�N���P �cU�В�;�k#=ｭ���k���\�BxL�l��D�l.L����4�b�42���k?qK�7�r�[J�z�d-P�,�Q��.W�/j�}T땵vz���|}1�fT��T��e[3���C���E��/jLxG�uϯ���sܒ}3a U|䑹�\NQ�Ą��W��wۜ�MA�e7ao���n�>RR�ۻc��\�����U�L�s��ϫ�o�z{U�d��0�8���"0F4��x�nY��+Ғ�Z�~V�;Z=��t���߯�<�h�G��w��I�B��a�5-�w�4��7ΐ�U֐դ������#�SN�#s�}����˱7���F�{�@6�u6�
)(�8� {su�������j�(ʘ�HE�~M�����Kn2�� 6��_��F�y�[���w��5�&��hE�.��;0.�`T�D�l_���w��E�wY��'eZC����!0�#y�\�e�r�y?_k��J�eB�����ҵV�왼.v{�P(��ge�������UCb����j��vuT���"sc�M9�ج%Zű���)yT��<И���"��Nr�ݷ��-ۖe�����x��~Ja���0�3A!�9�"L���]�	���M�X�_0�è:�g�:�!t�V-�b}LLȦ�:'�{גJ^��g�Cy$b��}5� �QR�+��g-��"嗖c"�[+z�e��32�1���%N�|؞�!����n���[tf�������MO�l������ޫ*(.~���}\���jR���_cf\[Ļ��/U:�5N8p����^9�-����'ja�6@�BV�^d^tK�Y���F�5'���fZ7�Ic��q�q�5>ٯ}e�)���&>Z��ٝ�W�����F�0��\\&b�]���i�MҰ1�*
O�Y�>p���+�A���}�s3��5���Z���Sk�����r0���� 9"?}N��N�����,�^�5����9��1��F䶩I[����ꝍF�4�v���آn��2�c��HW��F���R��9�{JY�T�9�\�4��A���+C[����au�]>��[� _�� �$ڜ�������Ro���Ow��h*�&̕��,��6gw��)"�(ْ4��=[����H:��W;�>I�zű+�����`��_\�G�sDS�KRV�����\�>�V2/*$��(�=��� ΗZ˗�.̍��*�J���O�=����Xf��Y7ˢ%�BPI9��9Qg�#�(��p��d'*��4������jiL��1AP4�e����0e1	DR�cZ3�7���<u�8�F���c{���E�H
�$���h �_�"tO��0Y��-����U+?]҃fK�$𗬑�Q/�*��E��\��Q��E-��=��4��23���]*�Y�N��
�h?r4�����k�֣'��͟K�i��?Z���wWP�B�1V7�rs��k���`���[�S��i��&�qż�$���,]@�/�ၢ�H;X��G��]ly��ʺ�;����3�	�˺���ҰElK�i�ʳD#V7o�9yR�"I����9׷�޼��WT��Ph��[F��2Wu�fm��^�g"��zV��ҡv�1��?w�O�����o�,�e�������I(5�Z%y��7 �=�!��eS��5Zh���j�}�=�.���hƈ8���VQf�����9�������o�$�Fe]�`˧{���|%�)��J����=���O�P(���0��o������rrS�3P�i������W�T��߃���s�|b�;>���q
�"I��AH7�y��{Ө&B(f�j�65�+��m��FJ;�V�h�{�_w_���P�JO��s>�����J���gs�^�݀>EN+�5J	���x��I�֮~c���=�����:�{���8gY+�rk�?_K��Es+먉��0�e�^����5W_9t��.�2�#��U���7j�כ���:�����J!�`�u�F�n���f�� �:�*���R d�d򫩭B�L(�Q���1>4�S�|rf���勓'cF+>��d��yY�:|@��� ����B�c��k��!����ym67��2Џu�?G�b�^;+ЈQ�.Dl��Z�$/T��&}.�߹nR)yύ�$zg"=���I��lI	?P���������e&��A}�O��p�Jm��½�sNէl\�ݝ�;�y�sm�T�vK��WZ�ձ�{w����lz4����@�<��۾��h��	^�\ُ}��U
S�2���z{�F=(:^6'����G�E��M��."@��e����&~����}�n�����)���GU�׽\�I��|$cF�JQ2�kײJ^�gչy}݂�Leŋ�Oɵ��rѐnQ��V�Soy���7���~U�=�eJ�+~~j���.���H���J /Տ�HO���j|�/%���L��=1o�B~�S������� �~�!zt|�f:�h��>��ѝ ף�Z����谽��w�H����� ��=�B�6��=+;��3���'�改>��f�3_���6d���5��]_��']o���VO�t����\��\�'zP߈+��@/���~�y�g��6gg˸d��w5�Dʽ�f�<�to]$���ԉj����J��9�p!�S��f�B��Q�q,=���{s�[g&�?^�,Gvi��ۡ��c+~7h�f3Ny�3uȆ��|^H)˩[	j����s�M��z�ͷ��Y��������ra�o����ݟk��f�<]���9���r�1*ͷ}'�練Eڷ��g��x��ُ��ú�%��t��li�s�d�ܻ�Xg8�\WNL��l$r*Ys��Q��3ޗ"�[��5����/�}q������-W�;\��TGP������{^����f���N,�8.��3<�|�o��?e���9��5ά��I.ioo�st��,W����V�b�W/����E�DtL���ψ��60<8gn�9��(��"	ȥڮcy�ݍ�2rm��Ui��ϭv�"��y4��X_*<��A��3�{Ҹ�8\Άn�E͑&o��hU+�\AoB��A3fh�0��%�S�*���7���#2̪��;�:I"2�?!��;���p�.�3�<{�w�G�H�;��0�?M^���jSۡU:y��j�T��W�r{���dNy�ud@��b�@1������Gv��mi�EƻN��{��Tjs`1���wW��7���t��^���,����K�w�f�_�̢x�D�m��_�q݃�ko�{�7��e6M�F�h��7��nv��"Ko[�5$��@�$C�ю&�z�tcN���X&���S2r"�D����hR�y�u�f�(�|}Ep]��.���^ޓ��.]?g�~�.E��m���k=�IQ�C���umϥ˺ћ���K�v��vwf"�ۄ
�-;:isNƼ�:���w�^S�l��Og��ƣ���ɺ2Z����ȕ�F}6y�\��e��CQ�;+�ݜ�0�l��Nt?��޻��gu��ro��,g��9^r^�^h+9�[v[��pD��Ѻ�n�%�����v^ت����s����m����];&=��.R%��m�vzu��ػ:N)ۣ�7<Nҍ�ۮۭ��y��Z�7��t]l���6x��n���#f#���=�`;Z����n�p������Ky�w��s�q<gQ��Xv[��]��:���;V�DY�R
��ݮ�����EH�3�d���V)d"�eϢٵ˷c[��kc��n��t t糡�����ϭ�қ�n��u�e���q/!���lI/�����.:ݵǱϝ���ζ�ɮ�dֻs��%�u۾л�/r�=C{f؏F�e��mV1�����Sq���Ů�T��Q7\��۬ �������[�n��i�e�'Tr��l�\n�v�+{0m�n�DS�a��'�x�.N����^ ��z�/U���4�g���ݳv�����l��k�6��8���4Gh2�ٶ�Y�`u���m��/\�mp6��(��h�;��x���L�x��6�݃��]�oX������/�I���pc�l��;u�����M.�ۮ*������a�����ӜWkS�q�kqh؝���jٓ���zZ�91�\��u��o+ka�v�\�&��ӎ�k�s��<�m���vw��Ϸ&��SuhV�z:�#�Om���E�C��aN�Qv�bn�ad��q�Ny!z[v��ig����5Ś����F�"�y-��\���%=�{�=mm��-n��g��Ƹ���e@��Gnx����nw0�v-�v8�n����ｻ]������uA�/d�Σ�3\�\F��R�sZ�29�!��&Z��W��D͸�_�$�w�U�>^��caUA��?`�T�X-c�y��?d� Z!�t��|�8��j9[������=0��1�	��9��d�7�z?��q���DFi��:/h���p&R��ӝ�t�C#PKY��Æ���X��Z���~3}8��"�9tN_~���5|�J���|��I�:;�f�浢.�f됌�� �l��CU��ǯ*I��)q�1�T$��X�y��q{���'9V�s�|e���Le�/�X1[�Ֆ+��Ⳉ>�f4Z��@�.��ݐ(^.s��k�&���i3iu�&(��t�������Nz�nk���tl���k�_˂��w�d�8f0ރ8-8aG����˅}�f��n��{�v탟c�8�w7P�u��9mVۘ�u�c!˲�\�Ƴnm"�4nvM��'3g<���q[]���=�]�tp���;��¬6��]s���m����P�6�ɔz�t����� �^��qyۛV�`몀9˘1BY�=�8����j㞦��cAn=��d�O�S81�x��:����`�D����[c���l��f�BNşQ����!
�a�:�Y8�'�]"	2N/#���@��Fm��FmRSҩ�!�QM��NzI�5U�A�~6�MmEV��[nA��;�\�L�y\{z�O������i�ݽ�����W|�c��Z���W����oWK�5��nt��F�o6��k>]\�ߑ���e H��YH
�h+��/}���~��ѻs�4a�b��5�g.�M��FR����l����{����k�!��	5�G
�ë,X�VE�O�I��o�o�o�5�"��- �Q�;�2�������L}FUk4v6� ?G�H�,�0�,�|�O��柕x�> ǭ��.|r|��:u`�.%3L�%�g�p5��W���{�ײ�����/7皦<�	 )>a
~,˓�l+Xesu����������{W?y��1�9�KQK��g'Ѓ!��;��~϶`��.5��}����1z�p�<��:����,���ۣ��.#�A���U�j�j���he{��������P���'�����/��Ӫ��6U<�cq� ��۫nѮ|vV<�d�ͻ��}���E]�m����S�3˻Yq��9F�W&[=�%t���O��~~��B��|I��x������f��/8ۈǓ_���sE��z2����}�V��{�Q���=7�v�'����� �&��l���up�9�蘩����2��.���sL#�*��B��$#m��o�O"1|��iZCH/j�!}z�Z��1d!���a��2b=;���u�@o(�|Y�o��&}!��M�c�>���xU�lkJ���^T^h�DUe��}�El�(���o����I����g3%9�4e:��!�����湗��8�/���=V��5Z%K�v#����s�~��ٜ�g�=H[h�(Yk^Ͼ����8�f*�y�N��P�����J~����d�~�u��ofE����z����}|S����^�ު�M����S�.��V������Q�T&�j�f���T������z`|�-�="�ż�T*�8�y\����\�ؽ��S��b�K�U��/>^�El��4�G�ٟG�q˪���"�y)�lq	ʋ �nZ!;v��=d斝�F����7j�z��i�r��Z�J�UIp��Q�M�o9o����q}�f�Y�_߲}x���>��G���͵�*�g^Gۇ������MY	]�^v|Ͼr,l%��f�y2>�._y3x?�Z���=���k~��xscMmS;&)���n�iA��آ<�U"���+�S}����ڮ(�������l�����t#�5x�
�$��}�������U�~����N~�����;�'�cſ�Wi���ٹ��n��vm�<�1&i����`]���4�kg)H��wx�/��S��ty�V�b~�ˈ��Bg�����t�`���Q-lm�%��9��������WzG���,�~�fk�սm���Y���~�`�J6?%5��s&����Q7��eg��f>tV�׍�2��	�T��s���$�`�/T:��q����$㚹P0zjQz�_U���W����Q�T9h����Ф��� ǌ�.����dV���v1]��v��8;���G�vcՀ�a�����$~�9�3}�Τ�q������}D������oWn<n��q�W.�oN��h�Fūё5O/�&���P�����������4G����k�%�>۟?!"�>�B>P��?3��>�h¼���]�zf�E!�SQ�V#���G�xH��p� �܈ZǯҴ�~����o%���E�z�ϠO����I�s��o�>�﫼v<d�C��vzX�~�K}g篱��3�q�y~��- m�-"	�}���Q����ei�a���rl��������?���ru�j:a�SR�{+O�̯ �r�J�d��
YU^������a���d�I�9�L����r3�Nx`�2�HO�w��ח0<G�Jڹ�}��>Ę��k��_�W��KЫ5ۧ}Y��Ff��s���FDMVkY���������7E��w�%D��1F�J=��^�Y��!��%�w6}�w�#�@���|�{k ���7.H�W����ky/)G�U���}��aG�%RZ�J�i���x<^�;?9��?��:������}��������Ϣ����";ף����W��5'�QM|&��ioe�7v�����U?(�Om/n��j���
k�α��L��^��^Ee�T�tv���3!K~U��G���ɻ��AQu�Q�R��m��'��*�#%@�N@��d85���>���wxr���j��2o4��ى��;t�\���e�:V\�^�uj�=��@+~�����>6���{������#1�֡`�Z���
/>�4�cE�hz �,0��X~Hz��$�Hyc�}k%f�J埲8�p�??N@7��\I���A!Y���l��_EE򫟟:��0�pف��і^�ﾃ�K�1��wymHyù�
�(�H�����-D�����nk ��0���bD��Y�>E�"��d���qz �"2�:�AB�D�r�#�#��r��R����ʀ���p2�{���}$�u"�a�H�+��0��v
����J�K�s�+����,��)�pmw 
�97~ۜ��)����L��3N�mQ���_OQ�"�-��'�����w�۰Ͱ�� t��.8�;�$�>n���@��2l���W��e�5�p��g-=n�\t읉s-�R��ֆ9F���;pv���\��E���m�~��u�9�r�^��TvMOv�}�u���Zخ�a+�\y�u����8s��L[��[��Gj,�ŨM�5�ӆ�Ow��ݳR� TƢ�m�E+��k�nv���>	&�G��O�����B":�]w�Mt��TVG]��`ț���Z��!�Q��d�m�E�+�
�pUH�����ƟڲR*!�E�.���y�{6�'����R|��O_���3�S�h�̂����ޜK�����΁)�����0�5w�:;�E&��ٯ�0r��<�.n����x~?9��r�&*4�bץ��"2IH�H٤����eо�$䍴>߾�v�ňᨦ*=uk��B,��^�"Y��p���ɯ)�����Tw���]�#*��^�P1CcK���,���"3YV�}�x���oGJ�A%)S�O�������9��s<�կ&�g�T����U�26�;���MXE!�`���^]�I(��z�B*Q�A�![�w�<T$+�������4������
�
pYв��|��Ӛ/O��l|C���ʨ��)�4K?x���v��R!ϩ�y=�j0񕬠��˂B�pSp��}�	m�K���:3��<�nU�������k��s#p��e�Ƙj��^�������N|�����;���L�ms� ��"������7���̀�̈́R��"�e9ʴ�۱�w
9pɅq��GǗ�/'�&C�,����J��TL�b��2nE����=vw�����o?����_E��UEm�Q��e.]sz�-����Xep���s:���_|q�B�� A�S]�oBX�#U�K^e �x�'��%�#	.<�y�yA��x%�&���=���B3��/�O��r�ȅԪ��mʦ��N߿c����⑓;�H�+�L��P��n{j#Z_}��H�d�z�}���o��3W��PlAp��Q&J^��=�1�S��{{k��v�>b6S�`R��H2I�z�6x��&[��&��l%i���uV��К�g�K�-���~�)�J�7ls"���"�yiooK]���iUrRu����UX��L�11�T����(8��~�������8M���v�ɳvF�tIh�n"qN�ƛ$����NQMa�n@�n;Wm�����������c3ִI!Z8Æ�g��4�9�t�91�Iڹ��`@'����-&v]/	�LLj>�d�l�����}���u��Q8��[�������>��csMOG؍���4~����8'���<8s�����ѳ�f	*s0ԃxZ;�@�bv�>c~�u]�y�#��t�	%b�������D_���>r1��F����Oj2Y���Ն�D�,����#螂%��˻ �V5[0�(Rϳ�םH��`�*B��A���]�m��n�M���2�oq|�RF��}1�|�-^u�7�ru�)�J����@�,��H�^�YH��m�P�����U���������Q��{�[iGF�vM
��jL��
�S��!x�����y�.
�i}���ݪL�#�x�i@9ߜ�U��w^�.�
n$��b� ��2�E�d�l ��>:��C����v��|3�<o9�1�I�	�K�Z LL����=��"o��ܩ����qmx���A[d)UV8Q	2���-ؤ���8]�1X(F�)1�~6)��<d)S���z�b��V릉�o�L5�e��	0U}>O�|X��P�P�־rxh�4_��.Z�'>%+R�b�b��?~=Yr�7y�G��I��T����}Ǖ�f�X#�|����$��S����݂��r�����#G׽}8n���Y����*�Ŕ�ЋC'A�g��X_L� �My�>��@�����c���**� �0_��(	P�d8D�[�:gª����e�lP�t�������Y>R{��c?s4��O4�dj�Q�����"E+�QA��A��ޢ��m��8|#E�3(�4st0�°�@�Á��a,e{�MA�������t�tG�{ϯ�i���9�));6v�G������>M&��;�7W���GX���K̷Q/_��hG�2ǉ��5</_"ڥ���@hmS�>��D5�ʪ1m�AFtǦ+c��)�}����|(0�?
a�a�����ͯ��{<�`�Mg%�h�����ɝ~�<�)����+�d��H!�x��cq�q[194�ӕ��BH��WZf�Vp��\4�8���f��}��ֱ6aAb��ba�;/%�F�X�5�����6$"�H	�ݢ(k�V��'i,�l�eq���X�����"@�$���o��`O�k==�f��"� �Gq&�	b��cS �y ����ڐh}Hwi��	����cf�*˶�3�����������m����*}�D�c|DՎ��Nů�-� ���V�!P"����M�����6�)$�YϷ������3{�UЊ~;,�v�|�Ђ�fȱG�.5�@ݎ�| P��B�����=V��pj�Fd0����+zfC�������B� ��GOG�d�g�d�Ϫ�O�pEP����~�H���PA�
Eb��2��)��뾽�{����a�}I��f���/�j+�5�W��m�џw7��=S ��m�o���O���X����/����~KK���#��;e,r�d�D�K��v�=���K�Ǟ�]�E�{��&v�=��h�����7d^�s���z���uϬgl�չ�k7!�b��DA��doie����2�0��9�o@.�ƴ�k�����c�k�ǩ�c�N�5�v� ��f���v�ڲ.C�熸���nv�1j����D��݀.`yl��K�j�`��n>�wt���z�m���@���"".{�c�!�u��m��o�ݞv�M�[��9�&x�Lr��F��2�)eN��o�ľ��\R��e!]�QI3�L��6�^��Ȳ}��m]-{�|����n:��oLQ]9�F-�c�(�2Ya��16oA0Iq�ߨ�7F�e/o�K_z�OM�[JYqؾ1��T&/�w�M�4\͍�'.`����x�Q}�sn�7+H;>� ��CD!�)Tok�O�Z�G�U֗�u}z�VX���ۇ�7���Q⭗���"~��*��P�,�!�6WD�"<Qm�T�
50��]��~�PϤ���W>�g5O�^�j�`����w`E^�g��<B��-i9�7"<9i)�yOː��Q�Z�o��ٞ�
��p�H�с��;��Zf��#�K�f���?yZ���Wg1YD���H��]:���ײ�k�i\`J�71�k��Θ�ێǶ�9gdF):��Xê9-�W��^������#�TEǥ�~j�%��8�� �Fd@���O���3<�d� >�g}Y�!{h������@��� vg��ͰQ�@��l��\I� ���s�7qI���
fN8r~b��+��r�u�n��Y����R�[��௞k����=Z�2�/�+ꌷoᆈi�$>>�ƶE�C��Y'Æ������H_}�0���^���XOdd;��}g~2���E��э��U�zJ���E��ĮЎ7fA�-zr�g����u��ά������Oo���n�bmv�(eg�@~�� �@��H��.�%�_zi@��:!�TSi|�����?�eq�N��,@��`����Ȁ@�'�H0�>�Ђ� ���s��5�)#莭rI�C�P0���\��jJ���M�R-�ɫƵ�B��	ޙY�_u�C^?h�!�,u��~�`/{�0]k�#k�4}8��޸i�r[1�U�)��RGB�oPQ����x��8綞���\lU�X�OӤZڻV'luВZ��C%&�w��Se���|��bBL$s��\��TK���.��㿝�7X�AU��rf��~��Zb��-�������HX6��s�^����Qdr9���9z��`�HS?_���H_����6!w��7�@��~�2#!_%��,��Zo����qwچ�%
��mEق��#:�W�]��Wz�Q1��}��WHڃ�2�c���YT��j�v�r���A�.����ͮ��Y���ѭ���%�An5��o)�k��*n���oÙ6�#�raLb�W����n`9n�g&j�Y�A�n,e_K۸j����s���	wm�$����o��\�}+���R�r��o9��+Y��s&��}q��A@��e@�YB���c0;t���r�(�C������[Ѳ�W�ko���{��B��u{9�/{������ݡ�-yFκ�
�dJT����k����;h\��~�w�7����xN�(EV�;��eѾ9ٍlނc�n-�{������7f� ��a�CF����!(�5�2j<���w��^��i����4C�_}#�֪(?�\�!���{�۳�6��L9eʓ6�[�}��6�0����� 괊o�
����V���y�Xn��/K���8�=ޓ�ٌ���X�8��M	��z��7rz�Z��e���t�#^F�.;��v]m�v68Gi�C�Ρ�]m�k��V��xA�ԟB�3j�-����>�N�/���k0��Z;��Y3�[Qm���1�X�x�ܔ�mX�mn9�����*�ͦ7��N�L�ޜʅ��;�ӽZDs�H�+���<���<��C�4��n��֍S7�m�������Ⱦ*�m鸹�9
]$W Φ��~"E��Wp����c����fM�u�Y�(+�ݗz0�Pn]�1�>�v�yM�hޏ=�N�.#�)�.��̑�dF�F�m���U8̣úo�\$/��m��OX��
�o�t�D���w�/M�~#0�9��;uzԗ;�ͬ���jf��<팭ٛ��]MUmb~�f
Ξ\�;f�ߞ\���S9se/}��2�oݻu�Z��3��z?���+{��m���k�Է��s��/�2F]G��>��:ق5���L�^���\tA"`��`��*ì2n��T�o�FSV�ݞ=Tb�V.��&1ys�B��Q��Gd��c�]}�v_{{v��|:H�c�nu���woyQ�E�x������B��H����1*]��>�{W]�+)lFb�;5�����Ms�0Fd���E
;ۭ�MN�S��Y[����b�:�;)=ȹ�b3dk��3-���bZ��G��}$*H���a�rE"�4e����bF*�`\!�34$ Cp 5K� ��P�ݣ�HA�� &�Aإ@ ���^m챝���X�l1|0�B�$��'-�'�7���B����·�ު�s{�D\=�ڙ��V���}�,��&c�A0�4}��b;���R��?T��SbL�_�$�1p'�`�_�y�a!4#�3ը�3�p~��}/dӳ�&����Fؕ畀��[�H��s��s0'<�ָ�ן�?w�C.�\�0pIZ�����'�j�4��K��F�ao����de�mW�T���o�
_�e�F�`�e	3�ȩ߃C`'KD�R��?D.��'�s$��9�:�*��U{����,TB )B��B�~��EQl��ךd�>@)������J����xg�5��˕#��U��3j�K�t��Ayo}}7i]��}�)�~�&�ld��4o�}B��|غ���Z��*�~}a�����^�/�c����^�־�{_�4���7�N�5l0���������l=V�M��(�;+�
�Ӿ?�>��&�9藩1�����zc�~�&�>��\6�|�|��~���񼷰�}1��Z�O��ǖ�q�6���O��	�0������Ϫ=������J5��o�-��PM|�W�yq��ґǀ��k*�C����_i�ز��"��vG���e�7ղ|� @>~y��ɣ����v(�)�x�G&�1�n�x����^iN{���ۙ�x�[�|���q������@����;�B����xNQ� �A�"��x�e&G��q��7Q�2R#���thr�"'t� �L*�����d4[n^i�ƶx�1�쳘Mi �õ�7���>c�Y��#o�XX5`I/@�@#V�y�'�:P����=�3��s��u���ݟ�'߰I��qեk����J�e#C(X�"X���<*�X3rG?X5���}g�/~Ǎ����SS��TH*2�
�����"8�m�c���{~�.gNc)�p7��A�=Aw^@��6��f���_e�u��D�"��'�**�⋫�K$����_E�>��EPp\& 8P�e�h
a���g��}B�
�-r#��352����J�	R�4 ,���B�A	�0a�(��CP���u=���%Uu7����5w�vν5|�vP�.V�;�9�cE�,�0�L�Ƚ��f��q��noVeab6�E�P��U�ۍ[�ѓ����pcGc�n��yy�W\P�j��F5lx7��痷�b&��gn�.ҕ`�qO<j���ع�.v������tnrZ���Y~�s]������wk�K�
9fv���bo���.�:��!�3��wl3ӯj�]���?ok��c&�ιM�s�̇Vs���?c�X���pgx��:� �$r*(�Q�7c�mAY��	u���wh��c�G�f�V��d�A'�s���.�L��TLV�*Y然�9Ԉ/�䧀�s�#$���`2���������GPlȀP���ϝP�2jF�#(qs�*�1?	бH�����^R�Wd5�A��ܐQ��oc>�q=�A_*�J!攂��;�S�I2#��}w�>�c��J g�+��������!9���wdV�>��@��b$��P˟�&���i運z�s�q�A*�u�	�Ks�CzӇse�*�U��-���>��sy��Ӌ��b�_�7䏤I]1c(���F1	����H��H_�ڝ�QL��{놠����;6�)�xKװ���8�z ����cD���:��ig��~���\=���YU�����kk ��@b��P|omJ���#��j��Ԟ��s�]GD����t�$�{%�%� /HB����#"�7��,,F��vW+�n�{K��;�nn'�y�\�V��R�W�ۏ��F�t��0�_w��~������ݟ����Ta!�ܱW㷛�'tB������`@E���C��c������~ףUlv�D�b.���¥��cS������	��5 c��]T�5�$)<�	}y�`����U�La�،�s9��;�D櫝�Nf�ε�ټ��=��3�ۖ>@���F��nf�3f��>�﷨�4ín\䭽�8��p���[�w��V@�| 50�˛u=����]���-~Fo^���.tLB �ް��a����ﴔ�,�����ϼXO�ً���a�(ld��,��Foޯy]���=��c����ݎ��e	�;l���">���-*�s�XS����И$��=C���%|>��C`bŠ�@,f���𗃔��uF��>����I�mF�Br���p�Y��1���}��'�@H`f�� ���������[Yk�Hܸk����ǻȤ���VԭP`V�$�%=Ty�+u]�<=t5&�c'[�Ud��◗9�s��ڈ�Wן�_�ɡt��k*mh���l��@a0��Dw��aV;>�\�ɣ�w�����Bj���w�k��⵰|{Mv�yK~��rb����h��znX(�B��3�#����"� V��~�U��2pt�;U__{������h��g˸�ߪ����߫y;48C�sS����ތ��a�,��3�mt&�eb���6΄�v��Ä]�Y������ca�f{�{����6܇��V�N�-�	��/[٘it�
C5 �WEx��D)!�숿�w(0�zz�qHCd!��M
-~�����XEQ�M���z�OY.	 +�C���F�F@�N���ɬ���!c����&�d�3��w�`��zD8V}խ�R ,-	[/��2~z�YW3�.��/��,Nٝ��395i�����+����������Dz&���L��1�Y�<�GU�A�#�%��%�Q�x[�h��9M{=�4s�c!H���Z��u�eN`��Z�.���C1�	�'�F���g�D	�2�Wmi����T�-Qo��I t7�}���O�t� ���P�J)1��߯h[K�Q���~��*&�1��Z:&���m�%��� �b�X�!�{ޯO��ہd_W��BZ��z��񿐾��ؽ�}��L��F8#K,D��B�k������ψ4:'hZ6 ���ox(�	$ɭ1�'5�%Y�TC��{�h�yA��LO��1uA�dM+㻽��L|�%�C;��3��a2�����������ߝ��;�{�}n�f���3��܈���wl�/>�T���5G��=���T)6c]�g���TVQ�/4���E�8�U���2�G�L���_�����kGlH��z��=uZZ]��>ro^����L+x�� �##=�֕��ˑ1�kwS�����<T�����'-��kꁂ�E�AքRL\�=�6D��t��a،���+�|p[X쎎�j,"�qgd.�k�74�;v�Lκ���=���uB3�VH�"O
a��Ul�`�������\�@ �_x�/	R#mW��5�|�47�ʨ����ﶅ��.~W�K�`A�&ډ��w�v��D8��ݳ�Z��è��ClO�sKX�6�(}�T��k.I,W�5��>v0/�~��𢮔��Bd����(���H�֦u4q�'n�� ����;�v��y�X����z�a�\r��7��� ��|�q�p�ad'���@���~����&&&R���,2�2�P]��s���Wǆ�I�=��I���3!�*k��g��ل�	@�6
Dzug���u�){�/؂�(h��ƴ}��!C���,j	A�V���y�@��>e
xm�=3��F��Ӽ.� {��>^�������q�6,��ϣ��N��{!��p�u�{:�ý�19�w����V=�c�x��l�.su�;u+�sc6/���n����;s�]�{���n�Q��x�Ѵ$=kF|z^��n������V��rw�٭��}��Uƹ�Qj�Jt��I�Ek�����nܪ�]���s<��F����z�säg"�"�띶$;/F�tZUs�����s{q�U��/&sn�y��h�,DT�,jAR�f{8��Nw+hD}�9���Ž_p���`�l�C��|��%��K\�U�f\��q�m���kk�\�<D�@+rt�A�_���;�UF+�2/{7��]ƶ�cҨ�R����`;���@���)��Pv���>�r;^����"F @ ��}j%��]�e�j�N����q��2Q0B���c_�1����|>��'��w0��ɘN�>x���H��e����Bp�*�i����!e�����frd]N�B{��}u��D{��5b�u�b[�]�UW����ӌG������͈- �������o���{?Fh�����(���bn�FB����T���p������{��Z���B�n�/�u�m��q�pɱBu���}k�}#{����(�����㾯�[^��l)�u�
��$�+><�rdG�X���� _Ӽ�?��ݸ����5ծѴ���{OM\mu�X�$�vҢ��
PO��E����p���znv��H�(]'�Ô>��HϾ����Oц�(~��}�;���/ߜ��\!�R�v z�r��y�ܫ�j���n��9Go{��㍕���Z�Y�v;f��]`���ˑ�㺸�ض����\��3j�r�k��Mت��JnO`���P����b�	���;;s�=��F\�MjJ0��N~�Z��>�)�]~��g�4�'�(�>><&A��C.��^��b4�2l$8�7�t8n	0[05f�	t�����s5�g�4~h�fL���U-V�m׾:x ip$<B��]	��He��b
���,�l�&M�VX̼�$%5.���Y��+E�&B�[� ]����|�p�F��-
�7��#A��c��������ղ��\u*c�}���U��taYd>����ͧ����ű�x�;^zI(J��n��4�"������fPak��;g�rCm;�7 ��"��+p�m�v7��4��v8L�K��p�n���a����JT�$�1 TA"@�܁����hIQLE��b��B�#Aբ{����%j���\�!�q�s��Xq,C�<foJk����ܾ��*:��:����	�`F�x��ŝ���=.:�g�Çԅԏ��rs�0ԸE/��*1}Ѝ,l٠�����Љ�Q:��"�_�Q~�KG�7�w4��"�L�x� k�_q��n���f���d%�E��k9��W��1��24��έ��勅v�D�P��j�����5W �����D�>��!������i�1[N�tG��
X�=oO�$d!>��L�� �p�۾5���~�8]�~�ܺ��@�#O���T.�'c�ra!&�^"�xȑT���k��#����]�Z�������9:�W^}���(50;v`!67e�qە9L%RI�[k�b���U|����]�|m���m�T��T~k���3��Z���z�, K�D�݇�i{�-�nm�f9Yc��Y�������v��]Z��B�x u�����<�a�8"p���_H�1HA0�<����J~�f���CO�)�.��
_A�Dx��������
cF�>�������.�Bok�>���W���D�"����EZ��G�t8� B���BΛ!��7]��\>��3�'W�F^u��.����0l�|L	2D7%�??'��%���;!ڸ~���h��f�2~�>��H,r�0,�+8�׷j������n���[l����>�>A�����x	�K��uƓ�7gg���M�,I��Pчۇ}���)�u�G�2��D��7)@��c���7���t$����,��^kH*�rps�jr�C�7�u��!���8%�օ�������p�ohR�m�k��p�$�^�*�d���x��	.u#8�P���	���j4|A��Ct'$�[��ow���� !'D	��W�W���$؃��^�B�kkG5�g~�SH��-n˫��xk=3��H	u�m��t�g��y/h-��o�������v���*"X#g�\
bDP%xlyaC=l0��Mf�.�S�Mo�}�}����A�#di
��&!��d��C��9��t\���UV����^I|y�`w�]| w��~��� q}��h'tlN}�~H����@����x���FK����(S0���������=+�-��З$Z!By;��XgH�}�hg��ݫX��>ǭ|���TI-$�m���#6u�;6;�5ϑ
�����@
~0�#���>��}�]�c}��:6c�\H�7�ty�����;���7-4""�$��Pctb��C=�bB/FF_ǟ|h҂{a��:��L�s\�w��}�Y���.JO=�d�hK�!��rC�8�H
�vod�<����jԺ��%��(/֪t����]14{����/%�&��N>�({�ާ�A�6��S�p��_v%'�����WV�k�6�4h�����Mғ:�[�]�57����
�0Y�4t�!M�=
��OL-:#h7[~4-�˓�+���F���j���b�qr�j��
K���kc���eLD����s�����K��o
O�ksgwZ�|�,�ݴ�wD.GUV��ꭾ���#n:��cέ�$us�9�jab|�QE���ɯ[qA���=�/2�zAy`���TkΪ�%�Mu�i�%ڴLH<a��͘�;�te�CO-�ú��\o(��L��^g�8��3%�e�+]U!���W#51�E�|]ۂ�{.>��:"&N]G��N���;�rwS�N��w`���1�6x�ދ0�b��Uc�����]26��7U-]�������7�UZ���S����ߴ�M�?V��R�Ʌ۝եf ���ٱ�ײnA�ᝩ��oƃ��$>|�?_Uu�`�������=�?��	�����t*�|0gt��n��[d��pb���wK6�����
����� ��Ծ#W��=�g\��uqًF��|�<�g�l�&ap��dTA�֩�R�u����$�����~�3�~��Olp�R��=D�=Юy�Gx��r��>�<�^m�%!zR�x���	5G%�m?�_Ƒ��WR�����a��z"�Ed���vr�T�P���}�=�}r�BWLVN&"���`ݺ[ew)0��-��Z�u�E%�����e��4Ӷ�wkt�+������k S�ڶ�Ǉ�&���[�[�>�8<l���fȾ����!5O>�ݜ�h��)��T怷7"��u�H)	Fw6��=���ր����Oh�6��d�N\kn-��e`m�NG�lY�m��M���wg����FɈ�]��k�x�q���]��=e]�;u��x��<��9�v���];eT#����;Z�Ŧݎx݇�'��Q�&��tn��콫��۞��ز1ʏ�#�K���q;b׵>m\v�{��H=��m烵�\N[�g7n`V]���9�z�gn��7]n��C���\�\l���o#��3���E���'��vݜ���oc�wOWp�@v��F�]m۝�+Ļ��^Ǹ-&��v'�6�9��)6��&�v�Ō�ѻ#����Xz,��Zx礳��	���3PeL�����to�ɽ/Gn�ٹ�����s�۬Lѵ�5��X鱮{;�v�۲�:�[E=�\^.�u��M�n��<T��1�\��٧����\5������@�ɵ�6�'m3�^͐�Q����i���� �r^M���Xu[#t:�"��֬���d�Q93�戚C�2��1�cݣ�\x�/N�W6pY�Anm�n]=g����U�]���`y`�1įF|���x�3�����XwEә��akm�l3�X�)giV.�-<	�K�
`gh:�V@���ф��ۜ���m�S���;�B��=�[z�yC�e�ܼv&w.n�7]�4��Sh���5�����G[d�>�t�;O<J�Ovڝ�i�)�G)����ִnNg��tXX�A�U��r�5;��Q}���խ1۞���O4'Fw%cHX'�s�/]�۰6��q������@!�k:���vk�����K�c����W+R <�ݖ��������]���]�D�4\v�A�ӄI$�9��nv]����"<�:s`8q�;�m��Y��+���=5x�4��g͈�"��(�K׿�/��$�\܊���h��0Q�˫3zG:��:3���*A ����;K _t���U�����}���Z*�*� U��%�M�ΨǚE�.��1S���V�H���p�'Uݔ�)���vt�f�J�;�jR�:WX�TXͮ�ѵ�ݯo nSiI�׊�]@���s#.g:D(K*DY3n+�F9s4"H�SS��9��S����:�Gg�I/c�~�!ͥ�/������Y}]�|�g�$�뇚k�p6���xkk5*��=S)�{��Bn*Ff�[;X�0C�qӋ2/Gq��T�nE�՛�)��w��E!IQ�۔�$nH]�:LU�:ԚF�r�~qN�������x9��岼)!�761�u�8:Nӓ���;I,"t�� 1�v8���sv��şlWV{z�ծ�cp�ݰ��6 �V�\']���Xպڇ��b�l���viS:�9�-ѳ�h���d�iD�J'[qr�C(y�.���3i���e9"�96yչ{e�{�,���[k���$�-ӳշ+����b`\Zf�p @&�I8�E>#�@�*RDR��ٛ��ϝ�Pwp�5�G}�Oi��`����I��kSl'g%���mu�rv�ny��/��V�����FQ~.7�U{_!�:C2z*2��!�U���5��g�٩��-B�L�����Vv$�)�D->Ǐ��4��O�kQ7x��r��Ĕ*���6�#�w��!�)�h���/,��sƃe����>~LM��#\�����t�	\3y"���I,�E���j/���;=��_���������}��+�A �u������У>���і-��k����:�-sV�S�Bd����R�n�Z���L�00�1Q���~���z�X�|7o �\}w�����WrP3�������o��}IT��jY��x�������M��1�\�f��{�0E�L|0�lZ#S8,�ɴ���>�[�~޻����~�����V5�q�A#��t��s��IŸ亞m�%r��������:��ev��W�Q7[�ޯ�����(�s����!���|ϰ_½𸾊��o��d����+7�xo�����f+;�9Nq11%2�"��ض4V1P��ЊB���ʠ�}	N��\���T] �NÊsuݞ��������@�{�:<�褝��UJ�1!���]���(��Y��N������hE�\�9����ɴ7����m�p�z�s��F��Z�0,�� C�2��3cĨH@�o�Y��8�w��q�P�f�A�0�d�$�L���`����b�^�]�20(��{I��ݸb=�K��~�3�0�@��"���@/�[m8p��EF�#i��|��˦�ώ��w?{��hB�"�� �g:QHP=��8`do����Tz"����.�hJ3��W��\Ji��U]԰bv�h��-�~����ט�EM;3���|������z����Hv�7��F�A�B�5,@ �A���%?���/�s����Ӟk��N,��%�:v�*YG����*�D���t1�ʥ
�Z^[���}�J���D��,lN��t��K�h��(�# �K����]ؾ��Ζ+�x����zX������
��PL"le�y��g��;�>��|������A�^m����!�[Q�V\e	W;�l�q�U�6�5ح�[f9d�3�C����n����Br�一�D��|&��#�ߪbUT����œ\�o��;~� �D�
�h��	�|^�t��@}���g�����4�溣�k!�/�A���2}��jZ]a���#��F�Qa\�}(:�!����`�AN���F���z�w�|��P��,!>�$��?-�N�W>��/����H�Z�p����1�������,Ux1��@6����v���z�hn�"P�a����c������/
&f�'�7�#�Ϲ�?��[ډ D�H����!��,ץD��� �@l��% �V��<S��;�f��~M˝n�'(��k��bt���'6Lc��WT�8� R�ciޮy����Ռ-MJ(�թ���Eg긁��*��ETH�7�H�>Ah@������ħ瀺��(�����E��r �E�n#|/�aj��m\�|jf��$^�e?r�H֮2�Y�Y&����c&	,<���_��C�J^~�z�����h�q��s�X-4Q1E҂HB�YZ$�0��'��{���D���Wgۖ��>�űi��ɹ�MNgh�zyu I
J�=C��vԎ;�c�Z��+�`Dt�/��L�՞��!^��.� m�:�s��}�7�A�N��p���]�9D祙`7��Yٍ�Ys;a�8&����H});:��쉷�/+v�2�䳜��>pI�Z�������k"FFQ�!2(�HkA�򯝟	r�����Y��B�>B��`/#�
9kv8�R)�1��%���P"�$e����&�N\I@c�Dx籉�t�R
�?�n�#ѵ�S8ʩޟ��pB��}O����T�v��7i�e�.����Lu��ˋ�=��j�� �����MH;��M���
B�$n��iD���bb>����<�:/�'\o�q���,@P����Ȉ��6VI�U��[b~���D�G�$�6G?��V��W�̺��*W�lY0>�e~��c�ԅ�f��\88�)����Z��Nl�J<k�EoN�3!������
~�C'�>��b��P���gƧ�O�(r??�fH�e�3�$�^yK//��8���/�7>A#w`n��}@p��[�b1z7�K���wѪfVO�>BD!&D!
�"�\�.2d ��pN��9?z�����G�ޟ��H��5�〸����
�l[�%���'s+qs�>��vy�?H�-GK��UӉ
�zdY�A��4xgE�[��S=�i�l�6���٥�}��ދگ�k*	��"�.m�^�U�g]�������c��;v^Ӹ)r�uQ���[e$�[��ې���u����v�E�����vݡ޽Q�R6�"�;8����h�/cg�܍d��P��vݶZ�r�G7��Z�u���,ԓ�F;J���gv�ٴ�Ŕl�ڮ�PmYǣ��(�&`��cA���aO\��<j��:#���l��y�mg������k�N��N�9��>&*DG�P��7m?�v��-�-�۞KT��I��?]��..Z�6�p���n�+��r�����Aڪ�h�Rj�ʙ��Qo���L��`��?l�����=�!ߵM��>?Vz{�XϏ�W�?��7[�&g���~�i�p�����'<�޾a����;梾�'!�E��{��A��$s+F�`��T~�Z���7�Oe���������g=�"��h���V�,�ُwZ{��	p�҅Y���&7��v���G��߲��`�-��대Jˠ�
lpUS�HL�כ)�p�W�H�.�QBo����#���>�l}�|@*@�X�y�F���.gw���������'�v��U|3�"D2�6`�z�[Q �N�t_���Ae@<@C���e�q՗�OӅ�ӻÛ�����4�Z�{�1n+o���ج�N�nc,��"�yC"!�y&�nۗ�G��B�Bv��(]�v�غ�&9�{)_Χ��](!��Ǵ���01cİ�g�к���'�$/}����x���#�}u?H��`@� ���Ug֡'	D2��J�x���Ę�A�
_������5Or\%f���� ��&4���*�bҗ�h99)���AKc=�E���C��ꓳ�}�g���</��$�F!Ы���,�(����x2#±���t��n������, �a�D�ޙ�F!�L��w�2Wp׷�X�z�kY�-]|#W}B*9��E���hG��ݿ��Ne��fS�ӣ�J=_��	CA�ܯ:����0���߿wЈ�IKE��[��Nߕwff�����~� ��yG�2$,��@��� I�?pAR瘧4Ċy��)����$K�9���^�b�(�m��ST�9���/����+��{xl��W��@5���ܣ�9�ؓ�I@:/xHM8d+���^fVrn�^��n�^ʎ8��gm��綖���n��ti6x���?��3���+X��������5�𾯌7���aw�D�%�?k��g?k[��A��	8!~s�����
�/�)�
�@
MJ"����~����2�ci^�c�~�\���q��у�9T����'��U{��
FQ��+�j�&��~`���|�{OgǛ�!	�r%L:r#o���Ƕ���а�@[VZή�{��,-��FE�uj&H�Ń���2_v��%j��������qp����|."�	��>�^&Ȣ/{�k�6����i�+�{\ڹ��K��1k�w�ּ/ޕ����Z2��A$�S�\�Xq}Z��DA�ތ���>�����4�#���L_�Ѥm�����$�n��������5?��I��& �z렍����a��q9]9��x]��r���;B=���>���L�/`e�W]����Wv�7d�PxӥeV�CXc2�8�p-ʝ�g\��
�:��i'8��+W%d�D~�q�h�w.�Iz�����)nSդ	���*bi_�E;���,3���قzC^Ę�K=s�/�8Q وiG��^=�mE|I~�����DF�Lk�~ϔ��z�r����vk�Mh́���蔛��:>���+���˾%���E]����-ukߐ��T�2����#S4n�l~"{�ś¾��d0Z���q&��G�J��O�Z0CI�0a�\"m|�gK������ܿ}��_�����#;昲��莈*�,��1�Ȼވ��7sg{'d����u9�b�R@	w��!�M/��\=��;��t�����dZ2z�^��[�P��&�.��p��Ɲk�Li}��[�8A4�R1.�Y�4��4u��dL�#"��e2b!��5~Ծ�^�#�681�v��2$��K�ܙ�c�` g�����#Wi���s���oWX��52�ŲL'�Ka�g��ې�1�9�Ӑ�Uם�=]:y����
����"�Э��M��٬�\$�.��ϭ*$[��e�{D;ܑ,K��i�����މz��@�J��ȱ��Z�m��Ԩɜ�m��{ɻ��>��]!h�o��x0��y�����xHr3����>��}8V���=�_��l��3�[\̬&,�}��L=����5!W��G�v���5�zMG� )�W����`�<�����},a���%4�L@h��MN�8=z}SM���=�Z` �A��g�悘��a�X]�@������{�9;�姟h�o�c��%�@	[iT2��L	?a&.����'���n������15� 0����3�IC��~�3�x�lY��d͊�OLɛ�.%�M�g~|8�(Q9���sx{ۋ�wq��Vi�'�Al��8�T1��������ή����ͦ�{S��F$5]˺S�L�����g׻+'OgS�`�7�8���:�͟%j9���×k��ڱ�s����8���cl�-nڝ���J)�rl��7\F�w^`�#�����>R�g�vL�ȓ�]r�[�����$&�!=�c��֮�v;Y5�s�ܐ���/j���᫭X�G=�l��}<[:�6�0�_Lk�A�Eu1t�ϗ��S^���Pc��.O�#L�#������n��ݔp�님��6�=v�v&r��q[D��L�n�Ll�{��ލ���wIc�Z^3{"�z�K��)�&�,^�1 Z�y��~��M�)���ߕ�Rw�o�	�b�0�$�f�xOw����;�Wש�h�!|�5�O�?O�L���5���p]3�/�3�JGD�斧�����B�B-u��#x�y�
�z0a&A�|3^���)�_\��}9�҅P#���"�)��+,U=�,�e�d��RH������jhϳ���<�œ+���ޫ�2�I��|I��o��{����g�n_����^����AL��6�{R����PO�u���SF�}�Ջ�#k<sɏ�Р�����a&����\
�(���F�L����U�8�l�QE��f���c��wF,�k[9�]�Ý�jH�<�'�җ܀��7J�{�������mG"���i|sH'�Dh"}���A����*s7~*���Vi�F��*�4�Sbx������a��G�U;�����E�������~��*8&;�P��я;x�N��KܐNکs+
��
���ѱ/q'5�U(��IL��}&�^�_����:ȼ�G��|K5]�$z��|�6�[����s�ˑ_ʊ��0W�A��3��{1���kϯ��d�����~PGBp��I/ �����HX��'�B�;�7���_����A�Il
�ɼ̂{����I�B��f��ݽ��������s}��PGq�~�H6�#T�}�RD��^���*3;�>d�}-3^���{�E��(�s�\x� ��Nz��3J�s����Њ^cC��W�$�����^?G�$_G�@�cG���Iv��*<�ޔ�0� /D/i�\qmz��ʏ��v����n[j�KZ1���[�ݒ��j�cZ]Yb��7�����܊~�7���?�X�?���[���>H�CH������7�6T7�$���c�%�3>�~g���v>�u�n�����Ԏ�Jx��ʅ��ﾜ"��a�����`J(�$I�>"!}�Ns��c���W�{c���>vg���"���1�20�N[�ͩ�7e�x{xm��ev�y�[���R����i�66�p�{᷂�z�l���IdZw����黇��7.D�l��ϸ�Ljj՝���^=�c��)6p��P�U�1��B�1���ES5#"GFꠍ@��<`� Qb���K��1�z��!�PS��4���ulI�"Sfmm"@dJ�b�R�HK9�[s�&���I���T��4�$�2�.��u��9>���T"� ���B�W���Ƒ5���z|�~�=ۯ)o�o�Wr,�h��˚'��M�+Tz�����u��ElE�U���\��>���Q���������*��ؾ��[|�,]J�%��]�6��k�{;��Kߧ(-��n���=:�N-�XX)�k�E<yxD���[��<gz��o4C�˘n����Eu,�3~%��ڳR6:�73X<��wy2u
z?�����-e��ѿ^�>m�B�gO��i«+	�{�݅�V���xb�Y����Gx��w{R&�Oo]��5|�eE��ܮ��)�*�d����N��b;t�f��;y��y3��'L�	��j����Ef}��ݔ�0�{�,�����/"�jc�'�����ʱ����	��Q�mP�����\m�8g��w\D�m]�;�h�Î�8��(��n��.P��>�=d�f��wdH��rgO�P|���I� ��w�f\�ܰ�V5Əgu2��ǭ�������n��|�k�؉]z��3v�fM���|(���SV����$��s\�y:�hi"Z�c�j�4��5Jh[\N�~kΐ�i�8�Z
�Z!Ey��'_&��W��O� 2$�i\���a�2�a���8łu��j*z���icA���	uj��xq��I���\+��4#�`������V���'��=ؗH%qI�t+��	���|�E+�H�ނA�=ҵy咙���"<7+����*�Y��l��Pu�TEm�F�E����7	(�AR��x��}yR����4���١P�UaǛ�;7�ʺ��,@��w�<�-1T�Rc{���ϴgj%Lѫ[9�r�vsD�k��5�1���2^�v�<v�A�ٕ����C���3�%�L�jgyN��me]��9t�t�u�ޤᩊ{��4���(�8�y9E�EGfL�~�yu��˨�*���\�v��`΁ց����A�J��j/;-͢��u��Ig ���r�P�+f�m�1%����ؚ�EB������6Q��;���,B�N�	�HԮkT�9��Q�/�{�غ���%�T/q�rv�nT{/�狾�^�B'�d>�y��U���𒈝���tL�HҩzA�O?i{1<��N�Y6�h�-�}���f��g\����U���<��?���_�# ޷���K�q�}W޾U �$��B��X�|�S�����T(��
�D�E��f�����De�s7-����PT��Lb+i��&�[�O�I~d�b~/{�Ɉ�����mQ�@�~,Ox�LV�b�ȹ���5uW#�L�$�*�h�	@M�.��}��Z�'<���3��o`|�W��C�Bk(��c��Y�~_��yֽu�W�! ���h�k�#�H�OM����<�c������%" 7�m��#�i�V2��dr9��jO��G|�c��ߐ!8�
G��(����X�Z��,V�`"d�\{��1{�hϵ���	lɎ�)�)d�[1�	��
� �(oi���\���
�����g=f�!��VX��&�J0Y��`RJ�a^&�m�8�����"O����}�K-w�2*�(G�A(��{��H�������K��ڈhތ�R�����i��>��w.blH9y�:�����uNr��/����휣�z�?�Z�2���Ϟ@g�#�}z�A4��Z��̀���s4���=U�j��k�K�U�<b���u~��{�}�M/}�8szɉĚL�����C�����s�xގ�"��\�\s����k�~���H5Vup���&-�n�vݻq�v�*�㓆�H��������"aR��W���)��IK�t ����
Z߾���jy�f&����W�l�ֵgW��1�w\��Ҕ�"��y��ir�~zk�^D�S|����`;1���7+�}_"L�����	�����wʟ�1w�򛝡_iB�˸4��4�-_ƴ܏���Ԏ����,e<����f����q~A�}l�	��.m��H��V���	@�����`t�or�JrH�f}�3���-�`�$��r$Ѭ)�v�Г9!�&��↽��I�Ƿ.rV;��'��-(��:0�݀�O1]���pT�G��?]W��@�����z��$��E�¶q,D6z�<�#��'���.qq��cs�c�zϝ�?�Z��{A�p�/�9}�q�[b��{�;�=����XK�R�OM�����vg@��Z,��w�{rK��d��<E�Hq��:��،)^}�=��-��M�\�Ӈ1��j�$q�;lgpv����h͕�p�.x$�-:6.C��z�'�n�,!��%��Ы웕8�Jl][m�nےun<��Z.ݴ��c�fBr�1����ɵ�5�����7a�!¦�ӱ�V�v��lT���xb��1B:�N�k�/}�!�l&�7.g�ת�U9;��?CZg�w��h��#�ϓ��2+HWUcj*� �s�f{b��6]����3�����������㾱iD�Q�o3ߋ����!���w�߶��<����oVX����$'�bo������Ɇ1���K^�X~��2&�>C�C���Չ��&B��W���(���E��!w=�5��cFPH�/� q��P&l%o�յ3{��@��s��t"�@��{���M�>����Ä�/����o�6�U��CNA��[t[��)}��B [J7l�,hM2D������=�O��d����~�L��D	x��VD�$|�gď��>�쓯�3}�χ������-_�\]T�ے�d�Dx�#7u��$0��&��q�͇����f���7�"P�����ExmHa�1�zW�0��u`,+��iȏ������$�6�c�v��F'; ���Y�����{6M�r�r$JK-i��U�ŭ����ebCD$���0��`��Ib�Z��<b(!΂I�
�����C-pqX�pco6����g����.���[�|��>Ɏ�Ru�w"�b�JΫ�Z�ֈ1z�e�5��,E-L�n�u�N����.�;���_M��--o�F��N���nUKu�����9����GG��9.�GרW�����>���"H�H}�3�B5ӟh��(B}v� k~�+�H;J��s����ŵ7��c�
6����$и�>�����"�/A6�&8�6(�,�p���WXw���fc.0��#Cf�>�z��p<�}3:Q>��.�`G�!����TA%\	r O��Do..T���w��q��3%-����)`	#!���x�Y����^2	d�{��x��Dͦ�y}�K�h�m��n�}�I��E/�m��g�|u�R|�01�aU2v=��Ű��i����d�#��f��4#�6ۑg�v]=����NF��_����%(x� v������`��Lo�LB�"��|A�!������qP3���;I�n*���=�!��^��(��X���>�1$ �4I�1q} �S�_j'���=�����{<��}��E9�V�s��)jdv�m�w>��@�ua��tiǁM�x��X�7qa�OΚ����y������T�A�v��B9d�xZ��o����VT*���^^4�����ʭ�=��AB����tŻ���!�Q�¬�6n��t�����rC2G�zI�����,$1�>Z8E����JX� �x�-������~坼0��(���o�,W�@���)�R�&��T{9ç;|,��\�7�ͣ�����dnY&b8��e�KK���3BGV�UEI��O�a)��C��O��, ��A%�xA"zM��O��>�UAA�Ք�O<���7	q�ױ�����v�v��Fn��C�t$���^q�qP�t�o���\�P��$��k�͙$��^�C>:$H���ء2�O��,?1%���:��U����+o�\����~��| c�����.��p�~��	$1�!z}[>��R,�������\/�����?>����S}��e��s�}������鿖�S�1a���SD�Y{_���}�b>^��*�\/���;謯]X��|D���
��2�7$�O1�~��,_���� c�^��랊������w�k�^�C�c���^���)�R*�v�R�[�w��vTd���!:�綯7U_*�xB��]
SN6���s3D������UZj�7�a$YYĎ#�&������7�|�۽J��(yw7�mZ2}�������oB��@q������zF�z�>�d���q�Α�
"��[�^��\!�ؙ�|$��HAf�E�>M���^�ԭ�d�Z��Y\���a+�p�8���q��m<�����ř���}�Ԙ����V!�����~WG�2��G��]ò�Y-��rwOx�~72h��!N�\���)��/@5�T2A���+O��QmGܸ��ϟ��υ�\�|�Ν�[Xo=�ʇ<�7{�><D��>d�y~�`z�q���:�?��'nN|\�ؒ7ZHz=|	~�,G��BL��n�b8H̩�|?w�~��huwW���"5�t�39������_��Y`�"a�X�Z3q[��]*��Լ���}C���>C�+���2 f NM��g=��o˼1՜h�2���?-z��G �
�E6��HM��V��i@Uw�{��@�j���dk$��0�KYرb��t̄���H��� }ВИ�A}�2��B4�=�Y��*��=��Z����L��1ݴ��W�d]��-���,�e�sg���q�	h(,(7nU�\]i�뒶,!����ud��0�H�ݪ7dNL�=����Ƿc��Y歭[����/�5��Y��:���ܶ�zn��3�s�:��u�88�{s�[���X���p��8.k����=g�]rō�D]�{=��<v2���+]�!��:�n:���w��ϓa���mý��.uF�Ws�n�g; s����ۖ�+�ޭ��\&�_��&���d�W7^���ն�G�/����ޝ���y��·Gk�f5�:<`��8��iki�l�9>7�ɨ@*�ұPuI&].4���f���m�0�^ML�I&|�y�ơq��U�t4OJ����cĥǽ#'&qF;��S�Q��(%)��lg�!ː&�G��*�̈́1�	_p3 !�ӥz�:7�����X-{�pM�;����	�RR
UJ���Y�D�/˜�K_}�H��� |T?v��/ѠW�Pfv��,^�I��l��45����+�y>���/�iq_�6됔�֟����!wܟ{ƴ�q��d��>�ǵ/gLN�ȯc����\���gt�ɍx{��ƶ�U�M]�f�e=s��Z0"��S[[�_�L^���%�QK�����W��Rq���'���Y�'�մK�����O~�o��@{�[>�m1$}��r�i泥�\5��ơ�#�#�xv}��["��u��O���;6��WMp���Z, X�z]M\\���>Mh��a����na�P��/�s��)�O�%�i��H0؞�j��˗=w��Z_��Z�����D�m�����c~N1� �&}�w��mb����:\?��Zt&�rE��m<�k�E���O�A7:�'[��{�zk6�����+�C~�g�N;j|)tE�5��.��׈қN����?$|�S��|3��i'���Hj��DǠ�O��W�9������A|4���Y����t�>�!��0���{D����X��}�9����/BC���X7P�Xu����\ĖY2��τ}��̢s�~�/ʈ,)^�����9��#�"i{�RK�`W�d-	?��#� �S�|g_�I�4��r��
�M=��VV#ߛw>[�D��u��kxm� �}��yd���(JA�5��7W�Hi���ʺ�T��s]��a��X�w�`�Q�HTޮ�N<Vn���Mky^�R�@�su�KpJ��j���+���f���\�������= ���Tł*\�"�{��b��}�ϵ��`��� ���Rc�CiZ��Y:��%b����3j���O�,P�ө~�֔�������g��}Ĉ��j��<� ����˽�%K�=̙>�çT��&ܮUD;Ss7�?h��_�g�y�>�A�+��!�;uӄm��N�n�����dm�Qs5�qn�/c7��"(��B���M޶Q_�C�@�ڍ�{x�t��Ҳa�A���N(�������fQ#�b�>��Z���sr*4���	�s�����e$��O���_��Coⵘ.%8 �$�/�6_��������.������*!VU���sT��WtJ9��_+>0��~>��A�==�'}w���L����������j�7��a"Ϗɩs=��(MOl��ï/�W;�,�|֒_�˞�Ϳ�'�yX�>���,�M��'��Ǣ�xȾ�OFCO䋏F��V��zxH���і���Ú��n'�nN�m~q}���lm��V�G&{;��_����߮E��i�>��h�"���y�_�Ffz2�*z��xy��}�מ+��5���^� [X?�z_e��ZI���p���!,?F�G��ޮ�^���,���Κ��z�5������d}��1��둓�[��@�87R4h���\���Y?n���	*Ҧ������}9=�v~��t�� >)z|��ٕ~�ώ+�ϵ���O��RA��H�}\ t�)G�U��~������n��_i��W�^�`$b������;JbcrS���2n܂no˴n(!� K��ڵ�D��8�s�}�n�C1�{-��{{1�u)������pP��[4p��0��P��D��!I%i��iD�z�ߴ��D ��16���j�/T裓��=��z~#?/���ʺ��u]e|D��	�O��U����z�x(�Hd��vb��g�w8i���?��&�P��nm����}�u��*��Jx�;���d�g�ɳ����HD*�%ͭ��qN'2��=f��aܙ�\��)>*����ɱ=R*���&F���O�鿐c�&?��Z�%��r��g&y4�#�]����W��~>�|���R��q��S�3���W9���-��\�E�y<<�������qVU���~^��яr��~�R�޿Er$Џl��8�i��������CW��/(�1�
��3��V>�0�m"�Q�s��=nk�D�|��A����0�s*��Ǜ��c^��O�Z���՝��]��`�T@'��q� �}�&1���̻2C�9_�ܳBn��n��į!mB��%׈X%�U�}�#T��Ǿ���;�j�z��{|ꏣ?Ѕ4�L7ryr��7o^���x5(t��ܑ����
N�W/gn��)R�:�����;�,�B�<�xIgO��qb�����ɩT��Q�)ʡ�g՚T�O@����nI�e��:��\�������� �'y:N�ܐ���'>�ϵ������^ Y�O$aN�k�h�C#O�߸�f:o2���3�Jz8Lo%��T��@ݣ5t��*z1QY>�~�u�p�ӑo�Ou|Ksd'qG�^��
G
���yw�W��]�G�78ke>�z�T��u&+�Z�uv�Od����F��S�[X���C��2k6�J霸��r"$��]�:�<=Y2�/bJK����{�c=����)��}3'b܍��,�Z���|�6㤇��ռrz�����+��0��!U���X�>�w?�歏�x�Z��j�`���Ҳ��[����&dlk�c��v^p�G:���5�k�֩lF�[�hWlJ��}�u)�1��z�$�8�22�h�b�PQ�r���1���G��I+�c&/��/���}�o��9a� ���&kNg�x	O4x��{|ھ:�3�ɭ����f�s�ϳo����~j�u<sQH)5q�(�3�#�G��><`���hcSݩ|��z���j����:C�(uJ4֑r<�x��֝��Nd{���Q���2|�5G��$C�I�:��o_Y�1�14����d� �Uy�Ɗ���]�8��m{4�V�-
� ���|g'�ed����no�\S�f�]�ٟ�4��s/���|9t���uA�Gn���6�J�v?���W��g0X���qs�^�@B9��&D�����=�<NF��.�����i��6���n�%;�����!�Q�N�]YxaH� �$I�]{��#�rD�M%hb._��rU&V�T^H���=g�k]V���J
��I���qb��,dE��	�c]�󂣞�t�5�we9�5�v�ڤ�Kkq�����Ϋ�tݙY����G��r�9�v��<q4Y뫴�<;�73m����n�-ۢMݙ���at.;��Z֑���{s�/4�O\n����lh�+r@�cp����z�ԑj�u��GP�R{�����vP�۠�r�Ĳ{�Ǭ�9�mh�^rB���&�OX.����\�y��6ι��#[i8Gp�v�U)q�j�4����s�'�곕е[�����]��Ǔ������5�=�vM�k�5�Ol˗<�<���y�W�B�ɣ�7X1[-no)s��v�H���n�;:������rk�� ��Ň�ں�c��%d8��x+nn��u��ƭ��f(Z�{v�己�\���svy��EM8z���h4b'�����Zewr&��zq�v{	[{��K�9֠��i��S�ӊ�������1�E��qm��Ѯ�cI��ֵȻ�n�#�o";�({[���g��������sؓ��ΓY�b�E�������#3W\wO9.gO�x�	P�!�"���7H�j��m�����M�<�8P���L*���E�D�s��a���㰘� ���j�X�bR�n{=	c��P���(탎0����8�:�+�����<s9�S��������(�pQ\R����������ɫx���y(����.�v6�Loh�6 �v�{w�۫��("���e��+���j���`;�v��Yݓϊ�8;��8��=�9�h�;�{W���pi�ͮ���8��2�g���x�n7 @٦�j:�{�.zc��avx�`��8�S�0�Ct��Y �\s�h��tq��$u�n�x��/Y�z7\o(۰��q�c������x��E��cZ��������mvݕN�v�&�]6`���kRR3@On'�qy��9X��Y�2�<!ŕS�v8��i;u�����vȝ���q�H��Y��K�罏�����݂vo.��S	_@�2d�k�u�VE�t�,�ۛs2�g��vz\[�#V���rs΍�=iy1	�a���Gg]H���K+`mv9�u����_N���m8��*H���^��J�!�c��E�������-�V讥o	0������}c�S}�s��;���̦KĚ�;W�ϵ�vM�:����\C���,ȍ�ڸ�=SJgL\�z�8�7�V<��G��@�'������I�O�۝������j1��F�����)���p�����Z�Q.�[]��ص&U��V]8��b�q��n�k��Ӄ�:���&�̙�P=ܳm�s�j�9�x��G���Wo�Ç;	<e4�7d�H�L��<WWZ�����qoUw���`�B�-�R��!"^�X]�p�X�3�rὮ�k�v�n���3���P]��;�=���c;j�eD4M[����ڹnǓ5��^z����C�gG7c�������k�)�������;�����Hz��#�>�=V�6�{3��۳�ͳ^I����\��/�*����۬�=�{y��y����R�)�p��܏0Ჺ���յ����<N�V�Y�lൕ������nNR:�u�-��z��v=���vۋ\C�á� ���E4�l���8l���_	�D��������U0���[��y�@�+���ǫ����ֹ�Jz�W���[=j�<���m{�{�в�W0��c�]�F��s�:���`��(E\�u=d|}�	�~>dF
�@9�5��^}���w>8�أ�!�졋�����`�L�0
L0n��M�2�>#e�ߘ�z_��g�Ҿ��NL�W�0,��$���&b�y }�Ȉi���Dף�s�L���RH$J�����@����	҄�������#���/^6f|�{�9�EԬ��}�����6����%XN�W{����F��p[^V`�ꌾʑ���O����!���_�:���{W?v%�0G�n` D!$���Έ�Bg�X��Ա=g�8넑7H�D� ����Y�m�R�M��$�&Q8I
�EQ&Y�-v*���ո8b	?6
3������W����i]��)2<�R��z�l>��Ǘ���O'{���E��r
aY�nx�U`�S���&?�_{�˾�{�N��i}퇔�7���#h�߲N��DE�+�vk������4��%n����k��]dj��z~v��?���������[*���_�� �q3"�	�g���������ǮA��Q�H������%�7Q���ʮ��H����t��PKs2�Iy���`_|�ehkg��+A�~��i�V�߻���ƞ 3|6����bD�Q�8���e�M��A���+Kq��|L�G;�~�r�	>�~j���u��%{R���\���R�"X�$������|¬����X9p� ����/SN�EJ"\	�������~��ߢ����R�Ǐ�{���HB}�ߺk�=V��ٕ��x]O�aV���s�}�Eyx�ܷ~����J�Ao���ݎz:ʓ��]���]�6���;Wmq6쎺�!�Єlv Ce����]��%���yr�,�L=S~FK1��w̓��80i�^c�#��}��7`ϐ����Ο/�Khʠ�D�:��o�G�"�W���G��4g���ׂ� ~�=r�"=_���ϸ�^�������CFq.�������g��}7'1�%�
@��q�3��^L��g���1�8��G��j��B�!�Gd�u����x�&aT��td�[ي�]�y8g:��&�$��_Z���v@-��;*`e�r�*y��������t_��Y9��N�-�#m2F8�.���[$h�D��<��`(zϯ�#��� ��r�,����s,�gϽNX��:���;�Z�;U���G"�KVa�i���4}�׾���g#�#����^�����	�����)*,o���������=Ӊ���0�<Nz��m`��hIs�����h�h�O~7|lh��d�1�ڏG���=��e}��鋒~�nP�M��ì���b�v֤�H��4�N��\j�uo[ݲ]�*n���S�yc��L���9]j��ŕV5T��\k��J�ך�Hi|������t?M|h?]V�/-������Z[�6�Œ�q���G�w���̱�~�j<k��?y�1A��'��||6�g����~����7�����<e+
M&a��ֿ9 ��q��p`X>��'��?t^1Z�}�����^��iF�ˏ~��'�ȵ��Epx�����Em�B+S[�|�˛K���}rw�D��W����m����>q����b��^��ok����OTSd�}�Vx�S�;�+��-
7�;��y�K���Yz��^���'��-��Q�y����{�#�m��:�ޯ�$?��B/�1AV�B-�WԂ���b>�o��ޚ�D�s�.���P�4�sB�\���e^̺�=�+�:�r�#>r�
A������l��bg��H%z3��D��\�W�#�ſ�s�y�|�.�N8�d���X:G%�u�d%.M�\�\7F�ݲs�JQ��Λ,Fw�㾟�)��0(2O�׫�9z��ȗ�~�Z�|)�g�=G�1{3��-�K��/]G+���ךz�������T�}^(�f9��d�+��V��L����J��	�^�_�#���� ����L��fT{�ё�dv��k��ן��NP�n�nL�1)�;2w�7�矗?��߯�{L}���o�{;�q�$����~���ӓ��Ϫ�''�{�NQ�ﻥ?ppZu�n��wua��ٗ���֎��>�*)�'8�Wܕ�V'��|w�|ueq/f��6k�x������/pd���?��@��&`��AF�ϳo=��˯ީƌ�8�\2��T�3*���_�y{����*Z�큳>;���7�a�����]O=q������{:��+A��+'�>�u����9�X��u_C����O
��ɩU�߼�ܫ����f}ᦾ�85��sG:��������lBr6*�)K���ƭ�W`
�aܘ-�"��w,Si��c��th2��^����x�W���β� ����絶�v�aK;��+ۜ%ݮ�v,�Z���z�v���S[��>mIN�<K�:���+g.�ݡ��*=m�m�>�u�c�7!#Ֆn��	����mv�u�1�q���On���D����هbZ�"���W.vJkS��e3%�-2��pGfN2U��K�Y����-���ꢵ�[��˷��5���1��PR]�7��iw�����מ错�6ߖ���V摳�e�o3sꙩ��Q��ށ�!yG�����h9�M��U�ݠ�B�cZ��Ϋ����4HO�u����X<4�f��>�O��n�#��|�1���k�{cаG�������}.b��j<�C�P�����|e^�1�m�a�<rk.����սf�/D�w��f�H�?;�}#g�Uk���9�M�v�ixc!`�����{D���F��v��� �������̒�� g�Ͼ�	�'�_�^gaI[�aElP^�	?1�}��z=�W��I*pe��e�r�j�W��f}�9�\yv;�/���Ė=������+��չ�k����=B�f��"fa��1b���z���f�h�.���n��<�@v��)nsܑ5M���;!.TT(�����
�W-��ϙL2����ǥ3��\��MN[�G���(���4�\�5�+�~��ec�-��������^�n��L}G�Z}](蟓�7�Q{�Ũ	P^�s�Vdϗ^�o�����˄]B�]W]�T������r͛�3�j��ض�1}�������$��}u�^^f��
I-<�w+Z�`�)ZC��\���4{.���^�-����?/b^4�|��z}�%4��:}�y�����y#������V�m?�{\���絶�ͭ��NdI~_yz�9g�d?��`d�E/9���fv�y���֫�@�^��û?OL�q�QB7�������W�ﵽ�x��{ǘ�c�j�϶���}z
�|A~Oۘz=����a��x� ��!�]q�?&2���oY2���3K���ޑ�����������7G�����5�p�	$=9�#����D_O���ղ���p�^=�}��ݰv42�4�q��k��=��	� ��Y��R2
��L��<�y�ַ������n�T&���R�r�~��Z������]'	R�M��9^Ϧ��	ߙ_{��WHJ�t??n�R׻�ۭ����a(���?gMk��U̙����?q}�h|���Ǟ��|��+����`��<���1ݨ�H|�{���[���d]G��c��%Bp�95����g:��ϔ�ށ�'g�=�|���? �����-���v����V�w���	�L<��o2�%$��q�]��b����:C��D���IQ���(5LH�{*
�q=h"Z��D�8B�2MG�\v�x���O�6�	<�_�}��l�f`Â�$A��>���������y�+ں��f���kew�5Ys�(j�*�x�h�٣q�D�_�Ψ"chp����S��W�i�
�O�|O�o	��d^ؓ`����Ic�����^��^��]׫���4��H}܉��v.�'ʭV���h��]�>m�h�Z3����V��Ю��tt'��k_?�$:�;�\^�ǖe�k���<KW�[����R���_]��	ί��y���{
�3��'�eO;�o��:X F�n̄R��������)$Ox�{��m�J%v2��M�_9����D�mA������	��1V��{�P0:|�x�O��v�1�Dzϰ����x�����c��~��=���5>�N�n7Y����0�����z.ߣ��'Tz���sz�6�z�;�Z���hDMOg�����Q������Z	Hy����P]^�a����f<~��v���ۜ�i|����C.���;B̈́ð������)^^�"�E�jk��I_�>b�mۉ��q6`[�b
���m�Oñ�,���`��A�ې�:����n�q���3��3�1�s�g�3���y=t���m�"�����}>0<ώ����#��Uf���|�!�\��2��w�vz_6h�A��Ul1^C�Tm>�g��`G��N1a.��70��Z����1ٴn
����1����Mx��{8֮�����Ɗ&U�齯�BI�-9I0���$�ѽJ7�^�߂Z����}���HHRbI��l^kZ�N
ު����?(G+(���
���/1�j/�~syő��>���g�v�O��D��>�!y���5���+ D��w5(~i������&%�͂������C͡�8��_UN?h��P���z�1�`�l�Z�ڐ��E��)}8a���I���fD�-���W�<��$�
�9
x��/���B+�'��~^hoV���e�C�X��[���|�Y�d̴�֞��0�%���[�'�L�ׁʊS4*>���2���^>�9MJ �[� �lF좂�R�!}���~Y�7�k�ej�7���7n��)��:0�oQ��u/�aݍ�p��o�N����~�ǋ��*��_�wc,�����7����qZ�6s
��x�o\wmkW=�8Wnx�\Cr3�����\�݀w���;Q�m��[�P����<m��j����G=`�l�g��xu֎�Z�N��|��e�el���(������{Zx�O�x]�0[��vE�O<�;.�[�6��w���N�������nȏ�y7/"�;e��m���g��9�G�Z�����ƒ�|�Y������g�lF�!Td���$��e��.0�L8%��y�H�d5�[��{s{�yn �r�%�X7#w߯������.ԙA	�!5���_c��uzz�	0.�^�� ���"p@��5c��_,9E��"��T|�.Ow�5,���A4�m;�M�E7pۗ�B�j�������>!�Ib'�ꭠ�
�^H����ح���yO�7HX� I\���_m}V�2W��l�^3�U���1vog
��}N��9S�<�L�8}�ea��I/��	"�Q��"� ^��u���Dl��""��{`cCs�dv	b����3u��ɮ��!$�!5������6�82�n��"���'��@ZI���]�G�����OY�<t����E�S�6n�|h��(�&7�삠laH.��֓��?���ؑ��N��:������we.4����n����`��*���ߖ�S�7�%(�@(�(H���Q��	ON�p��F[뭢'ː��Ɋ����8��̾�o^�χ�Ј�W}�h�~5��~�=����̗�fH+�r�J��}�k"�97�`|>0;��rN2!8�
��$Z��u�#��[�N�b�.q�5�f����C����������3=z���#終���*�͙ ��w��u���	bTD܅?-�7�q��}j�����!xv�}*A}�7H3Ol�nI4.z~���@t��:�\{X5�<���~mT\O��Mw#}޴���y��aS���/]��A��g�Wf���ށ�TC���ޅ
�(��Ud섒�.2��> ���ϫ�Gx���ߪ��s��Ō�_P�p�f!@@�j[�y�#���A�������Xw�nz*�u��4(�׎�i�h������T�eZ��vo��3õU��0�m��}!����W�띭��q<T+0r�Rg�����[$vP!$��pRH	�pe�d�2}K�$�Nho��A԰R'!
�劣�NJLJ
�c��?���������)����ț'ᵐ}\5	�!P i���pI�9�@ۤ�����^M��.���?:�Z;�u�ݑ�5^�C�e�Aw��js*Ej1���9_�nWl��64u��)ˬ�TtTVm^�)nRP�7tEAs���^�s�o��U�{���5]��4dX�< ��o�˂�:����}d7��y�1��&��b��>}���عRӑxv��xF�1k�_&�[U[F��6�:}FX����Q��a��jѬ��pn�<�1� �w�Sh+�/�O�]�l�[+s]2/iE%��P�3���&��d�p�����;�e�s{'�����Ⱦ�I��=��ߌ�wi����/.v��{0���!yA�c�ʡ�I��� ��?�6}��;I���s֦c���Er���x+�WE]s��|T��d m�2�9��$b�X�ʞ#Ob�峓]�9H}�Ѩ�yG�`=z�NqˍDΠ��r�EɁ��:׾��^��4gТ�m�h���	��#��7�.ܪ�ÝɕG�:ջ3�������s�N�6s�1��P�ay9Ysa{KK!䳚�V�������l������/9dUm�x�Ջ�N������Vs���2�sq��>�廋I����[�ɡx{v���FΩp.���l;ܽJ�6ݲ���:|q�Rxz�,WF�Z��e:����7��l3���}��Y�}ӷ����צ�ô+���}��=�r������k�Z�z�v�gՕ�v'w
�˻��5��-Q��V�z�M�N�-7v\�;B�6�i��C�n�F�&��=t��ɽ�#M�t��Z]][�3~n�l����|}�����:sj{��'�\�7�[}�A anD)5kݙ����Vwj,��V�%z��f�\���7P���֮��8x�ć�2�Et�������U#�i��a]=���l#��:\�aϻ��f��͉M����
�x�e�ES �!�����#�͜L�0��<p.R�u*���T1��V�,�����#w�����1u�5p����jSɹ��:>���1�w���A�2����mY�/fݴki�ctc��<�>����������!ˍ��M9\}��l���^��2:��Si�e[�l�m�wx�ה>�Xpb�\�Q�Ƚ3������T	�y�b�E�Y��,�0��Q���WJҏ�٦,���6r;c���-�T@�zc�p�[>�h�� ��e�SP̢>�H;{B#9ֲs��=ѷyP8�O�94+���<�B��8�Q��w�9��wٱ �,�s�L"Q�3��M}����gd�)�!%���>+��9Ebm��q��bt#��+չ�b�ĉ��R$��&,6��w�+D���Y_{�/��׌(p�m@i����|u��Y�0�)���Y��$W���D�tK�y���}��"/�Lo_;Ϸ�'s��
��-�B%�d�n�hg'���㵷n9�͌EDRJ�k����b�Z֔nh�Q���Yv���@+�����������}?R�{�{�ˏ\��6��c3��/��KSC�ʾ�u_���s�8.V�ۯ�#>rm�����"��g�"~�nE�m�?{�t�V�}��XPi��A�H�ɯ\����3X��R�\�q�n�^'�#@��w,�>�_7"ض��o�hPen
BFђn%�?&N�s]�gE�+�dG ~!|�ؚ ���
���D�u���.�VƟ��Z�}�Ҩ�>�F|�ő�ꃧ�ơ4��֫�q�O�q�Ќ���9��t�`G�&lDy�dQ�"��	�8��6�B*�#��-"QA;��E�a�!����(�'=ę�~�uwA.=�>��^�c��w�ODNx�`��_g��zu���~���%s�hwK�����'��+��h�cH��k�֓a*P=��z�
DQء^8�뜟~� I���{��ޕ�?�;:��ꤳ<������4	&U��#VZF�@h���F���\�{�k���k/}gv�Ns�����l��<~�yB/��}ޚ�2�+�Fl��4F_<=�C�ʈP�,DϘ��x�|P�X���&5��"������d��c/hN��7b{w�_
֑��JJ&\
^:��3.WI9�s=5�V�~?h�8kߌRs��w���/)��g��o����E�X��yō�Q{��~D�չ��*x�M���[�p�����+�'���6�v�1�����s;�PYqHŮ�Za�)��|������z̺mXX��ߒ�;��F��b/"	�Dd9A�F�֭����-��IZ�Vܪ趨I@�^H�7,8��co��9y獸��qq�j}6���FǛV��q>X�tZ��j:��n/=��k�ۖ
מ��q�t��-�=#Κ��$ 銹�HI����Ӈ��k��-d��8;QG8�Y$]�ϖ�6�Kf����������6{\۰�m<��9�=�R�Ј�R^%�h׉���:�h��48L/�����>�We�9R؆�:g�+�4��i��6��H�a��Z�'n�.���dl=��֗�׶\��H�~��A�0���di�>^W��ܘk��[�2R�zs�Mp1LKyW���>=�4X��+�f�0���A@�w_q�}��K?^�X#����q�|X?+�D����X���FB�?`�>���=��D���{򞵤�ܸ��}��qqA$�Uu�O��{�X	��h���h�}������y{]�ջA�UX(�t?e�o�=�w�}S����C��W��7����k�Mw�	ʼ����ͯ���i���B6lOL�=B�n-@#=Yz#M�^����q6%M��f�E1g��)	�ɡ�}]b��9��|���}���S�W,6�(d��&3���@
bC{m\�&;S[~��M[����l-qǧ� u�����*�#x�BB��8�x��@�f�E�_��6�̔�M��&I"u�?5�.�3'z�3�U���	D�W"1��lW83���d�T����F�U����&�vT+q����}���8{f����Մ�Ƅ�R���g��-��C�6r���\]Ϯ�g�ݓ��w���2�k�}��)��IK"�W�l�|����?���z� ��4��V�F�G��v.�o
�����C�Z�'y	�ǘ�A�����F�睍���M1z��ߖ������� ���!!�9�t��	��;%��BR����|����k�^;��V�i0Q$
r+H�{�HH�N�}�b؟O	;��������>~@:_/㺒9O�޽7�$$W.F�tpr�q[�
L<^\�v��"X𢵂j��ƌ�e�o��֦��6a�J!⹱~ω2E1x��_��k�DPuw�Z'��3��.�(Y��@tF��;BSQ	[0��p�e߇�\Q$vGζb2��3�	Ϯա5~����|�9����]�V��}�k{�;^�TQY퍩�/�^�'�i�^����5U�㠙����	c1a3���V���[�Af�*�R�k��/7��Up2���{vX_�}�ƺqC
���8 ��,�Y~GJM�8d��X�X!���>��xwm��p���
$���}�1M��~�����NU�����x>���M��4+�yT�c뚩�=B�~�����b4E�*vD��������<C.��ַ����WV�cm���y5�d(��o��l��w&��O��$�`��
"��N�9�k�f1�'ѻ{"��]fwB�띛<���Y��j}� ��:Z:�>���~���숌�}�D�f"a�}V_�9��߳��J�9��F)��. �3�)A ����*��g��Z_�j�<���:��7��&�c�j�{�(
\0��}#5U\�|P�|G6JD�^�̈́R�8�z����h��E�ӻȗ3���k�V��:�ٟWyE[���L">+��[��Oxߙ��r-OH����*&�״��HF����&����:��HS�ߍ���ş)h���=������.Qh�Z��/��k٧�`��7��qQ�<ZB2�=3��YF�o�U,�~p�+6���h�Y�Z��S
�w��ʟ������}����;t�
���g�#o�{P]�=}�.��q�|�RYY����D�oDo���E5�E=���r/�l��"J&T�,h����f�nӡ�FuS�"�s$�u��a+��48Ҕ2�Y�@Q��klvb�6��|�#t?�9�7�_#�p��лi�`P|���\�P��pON~�ݾO���ꈵ4��U�~%��d$���!��Đ+隞�P0�u��/@�;'���A� ����]�x�U;�	lzw�R$��#:kǽg�0�<lE�(BA��]�_}�o�Fڲ�0��W����s't��?�Xai'���|��6�D����}��?O��J)�k��uWR�,�-�
 ��@��Rh�_{�q~�86�Hд��ۋ�`n�Qx����>=��=PF$�c���:��ԧ���k�(!؜,5�sK�X;��c���?��<��?^��^]]���5Z6jX(�e�����/]OO��\�L��RY��Wv�2��n���V�]XN�pp�t�^�.Mf��Q��v���	`�j�v{[u���>�U�Pn��Ln�"&]�A��c=�=q�ɽp�s�1�I��n3�l*�`Y��x���{=c�ۍ��;Q�I3���N���˲�m��gg-��ǎ�����R�n���Z3Y������[luGN�=kd?��̷:f�R�Ǣՙ5Q����(Iu�����B��쏋����D�1�޵.�eNLg�v��:ꭈ��e�YmM6��ִ-'n�u��ϕ��韻��tVs�C���7��X�:f���̱Z8�ژ/|߾dT�T�����%9�7Ʊ�_ّ���AV��{�������_�g�{\�}���I�y���MTaBLxȕ���	Ж�:�/�Et��7��~/+�g�߆�F�:���������2��Qȿd�ӕ�P]t�w'Q$|�	>lcl���h��[�;�Y�[t�>z=;>�g�����2���J�#�27���k��4�d�~�?��?Y�� �9��Cqt�兄p1+��R%���=�Ap�z�#�)lZ5.(����MҰ�<X���e�g��G�l���KalWn�#K��>��HG�t�C��$B�g�`�N���{"iq~��gg�zHk��󥊺� �{����i��cS�_U���C��Yw5N�k*ij�6��ڮ�����]�$D�/)�x�M��s�.p7@����su|bX�/R�o��]����+^�~H�!�u$��nd�na�6��V�%������Dt?v�E�{m������\���x������-bx^e��G����8*��Nd����:�'����-��թ�zI�Eￚ���4E�;���ze�b�E��>��7O��3<��I��P�������~�y[i��*>���t��D	g���IYR�u_��V���՘�P�{�#[�Y��='l$���]������%���g�併]1��R	�2�7rGG&k�U;d�L�����v��Ŏ2+۩�0��ɩ����B8p�P�Ԭrk��k=�f����з�~<(*��ևM|v�̛��$�B�}�Ȇ�l��$��&I��n������L�@�H)"T#�v9\K˽i��)�m^u~ }��n�p�0 �2�'��{��ƿz�%�d6�wV�Q۪��/��s�w����c���T�����+��P��v[��|��%�[f��0�y��fMF,����n%�C�,E��4E�n^݊���J~^����k΋Ꮩ����q{��vB�u�75z/�nY��Aɽ����V�%W��4"~�("|+B}��C���V���^�W�уCqM��!2M}ChX����	������E�l��z~ڲ3�?V��<>�o�?WT��C��4�%8H$@���h�"��܉���s`U"���
�ɂ��֍75�r��7��*ʒ�|<�y�T�3�����*x��}���v0ik��%$�7�uU��w���1JW%m���[�^���]n���|�O�,L���H����<��ᳺ�*���N�f�9E����nT˔�2�i~�4�����\�
��������]��h5!���J�D�QȖ���V�������  ),q�	�e+��8T�����	v\Z8w�����w�6�D�:;w?�c����f�Dn��h]��mq�7S��d�g�WZ�M퇮�O1��<&�]@ڈ��1�8!*Fo��g�H��͏G�L�gp�0>Y��8������"���{�.�����O{��<A?x��LN��LV�'�;�G�o�gy9"��ü�f�+������ۣ�m��%��0OO��݇&�<ݺA�[�$���]W����7��2�4�bȣ�%x�>�饐����}�y����7��Ə���_��}�s����7EU�D� �4 4;ӣ=���J_2�f�w;0���bLkc�Wh6��o��r ��W(=�	�3aя6��������˻܋���=�����'��[B._۷�N2F�#}[����٫ey��(ɬı�a�pKh����Dĝ����<X�3\�~7�9/�$�>������E�xQ#>�,��J�`�޾~�薹��Ƚ����BLvI����|E�?��	������������:N��T1�03`����ϊS>Y}�q@]7ʴ���(��#��bx�ֽ�^H���sn�&)`�ov)�(8ot�����v�6T���:]$�X7��x5o]��瘄�̈�!��M��p���&Lٝ����S�['���U�#[��Sw8g�a6�Z��OO������v��u-��[�A�z'Ϣ�0S8�a�G�T�������X���a\ҝ�6�%I�b�=餦�i��L�E`�a^���ʜ�Vz1�s��<p�6K�.Mv�>�>�PRXtr�%���<A���k1N�s¶���ק���-��fvv�$�[�=�����ci�/�9��r�w/W��	���c��qb##���)���;�gR2s�W��s��S�|X��ʇgl�[Yfy-�����}g���[ا9�e�[�M�o��\Q����=���jy�-��_)��m�h䋑��Z��!�l��{UP�y �^5�7�F���Oz�n������*���5��8"�-�%����I��[0����B����El	���m�Z��!��u�h����o���������46�(1�qᤧJ�t'`ML��̴�S�Ʉ��[�C�wOO�v�Lܘ[7`� ���ʶ5�c����^�븯�/ynNn������ӹCy�����;��P��^�a��z����(��R�gxm}�}�����N|��5�ʄa�Z2eh��2����6�N\n��C��:sX�d�1�M5$<	mmSl�I��u�\��O��اa:�v�7Jc�s<��SBi��\`�D�fRZ�P�5<-k����m=�[���1�e����GMŅ���K�w>:�w��5�j�a�����$�m�=�1os����3:+�ڃ/�
8�)������2g��.��t��#�	5�뇶4�������Vb�۝�H��絶s��$Ƕ1����{u��`�63ܾ���tt�Ӟ�{m�S�b�1+מ�+B�[t6�ý���[n�1�=�6��&��ݎv���o�n��;Wd[��؃���t;.�q��ͺ�iӌ<tZ�:�Eŗ��e4����$:B�s
�5�9�����d{IZ�:�G`��NҜ��[s��ޟ�!]�n(;���r�7SGw%�A�=�/d;<��u���+�/�a�^8�Î��͞��]�tc������3����r�� 2����0���(�,��H�P(�盶�p^Ѭ#҇ez6�n.��W��.Wlu'F���6�׮g�4�nv%6ٹ�\�H�K�����)��َ[���ζ�n�+�:�wmp�a������-��vY�=x�zbD�t6''�$�f���ct�y��y����vӛnܫ�a�tg9d��3��wG&>���(��:U�P�#>.ǩ����� �k��t[�@�ts�W;�}1�໒�Ɖbղ
�hi��R��`n��x]�>m��|�Yխ��I��/&{e�����nGڈ퇏<����Yˌg<����vȇ�3tv5=��<�Z�n��g����1Z�w9�fV2H��]8�{a�2�{v!mksn:�>��Xڎ�]��؂�r;n`��1��5���]P�Ж�2��=��<��֞΀�Zy�=v@�kJh�n�rW��w;l��uS�#�v:�K�Y���W�݃��u�D�k��s=�kr�gً�s��\E8*1
nÌ�n^��v]�ct���u�`��s/�����t75BȘs�"?�]��Z���yD��}����8}�g��d:��ϯ�!��`��pnO��'a����U�N��@�tT�ǯf�S�o�.�_�L���G'X�B,_uv�p�knN�o)<�����$%��������Y�EX��H�8��"cPW�'���00�'*aDY"�pB��f��S�2رT�GkvD�݁���D���5�pj�H⴯9�;��_]G^�c9z®�XFB��=��7�+6}KEle���#�%m����yS���I�U<6oMd��;0��{k	��Z.�"w�Z�����7Y��q�=|�>Ƚ��u���U�#����~#���P�R��|d �:`�6�����\nps��Ze��q�@��uҸ�/p����mv�ݔ���ݰǍ�;g�:]�i;tvEx�¯��=�`��k;�֣B�'X��۲=V9�ݶ�p`�:׸��r��y]9��:�+�X�c��)���]�!�rrrq����7��Ծ�G����qv���s�s��˅V�vz���F���������<<�ק �QǪ����v\�xq|qn�>2b�n���7b����#N��ӀD7k����93"�ݚ8+U[&�i�F�m���N�.�����ִ��U@!]�/�������s�@�\	���>��M|i�x[`�#)���s!�uS��>�S8p�D�Ќ|3c�A�������S��U�E5A����`�O�x~6����WΣþ@YO�LOY����p�!�f���h���>[~�Ϗ,�X�+��x�_�����n?a�<���am�27�L6�8���;����|�䀼g��BH �ts���I_|�o���#��|)5�A�R�ᙙ��J��= ����6~��(�����[�ϴ�{Ѿ���AH��s��P�®O2���N9bB	c��@�L�ޓ�x���5�>{no���w�'��&v��쯿DH?q%{b�����?�.��;G����>����~��b�'���M$C��q�>.�R*�����#�&���o��ʾnK���#�ڼ�܃�RD��,��l�%����gK׷�ϯ�m9��c9�1[��_�Z"�n�џ.���""��s���!��5,ޛ��J�>]��ϝ׊�C���w��2�z���Y_{�
���l8iC���[ߞ�fP7[�`��EF��]����b��ڹ��fY4E�<�'힝w$vI#e����7��s��������?LIz(�׾����s�fx�?f��ka*�O<�cb��m��3D�b�Dx�}���$��w�u5�����3�~}�3���9��D#s �ٵ�M�k�-�ASv�c�F��=t�:�lu˞��`
z��#�8�}�-���B��uZd&H����Z�<5��?�k����:Qτ�L�Fo�`,b��P���%ģ%]���N��Ϻ���������6Q��o��/p!x�� 8����$��^E/����-b��7��10&B����D���s�!"8��$�n- =	���=��s�N��?Gǯ���Kb�(�ɯu�iGgE�ոnf���1��=�at�Q��NVt�͑�������-��A�R��װ3[��R�3>�������S�~>H��}\)r&~�X�鶧4��
 +��&F�����E��}�/_�s�^�ykᑙ{<R���_ �Ot���~�����RH1�ׇm���w���.L�{��R��s�w|H�~ź�~� �P��=����ٱ�g��e���*��� g�Nu�>^;��kH�uJՍ��ޮ7������YQe)�S�}��?gU�e]��)蜐F��
|V8������c���uy����Q-��A��%^��Toٿ;�v�P��qv�A��(!�H�j`�ğu?�u��o��j-��D}�M:�A�� �	�O��ފ�ֆ���ļ+;!��@1�g�P��gǆ)��w~}o���=�����z� C��l�_��^��1'W�/Їw'�Z�$|f�oި������e��Oo� 5������Z�svG,8+�D`-)�7�і7`:6L�D����q��-c�+��SG�\��J�l��J��jD��x�M?�k�Q*�e����k���=I�:��m�/`VMɫS�� C�H����� &+c�)q�n9�?|���uq�<d_؇�YU���
w���To��	U~���^.�����1z��+X��-uZ����c�[D�8��1%�İ{A��Z����޿�B��&S,�p�\%��}�׍�7���x�9$HӺ�6]_�~��yoV��n�'�w����[���D�+���D���g����H�b��N�������������"r}d���""�H2)�_|8������qΧ��w�eF�G��^5�ci"��X��i���n�)[y۵�9��D��`�I��r�_���`�(���#=>�[�EF�$����n�|�\�8j!�Ӄ��Ҽ�N���1�%��E�4@�$���u����9�G��df��g.,�^���SQ<�$��6���1����2�3?�.��3���?=�.I�n>�z����ǫ�-�W��s����S��:s]�h5�Q\����#%\q&����p�AӖ�l�	�<[#r���\����c\f�ϥ���3m�:�Bm�m��-v<�,%��`���vŷ<����v6��I��i�Z��Qֺ.wG<X!OY��ܜ%��!]u���Lh��F�lXC��C�2X�bm�4�H(���u5�V�3ʹG�����є�d�Γ�6ݮ�ٴ)��>�
���s��=K8�P*e����Cr�m�Tf6;vv�� >3Ѯ�P�:�����}�=(&
q	��)�{�N����H��$�{%�빟�B4�����A$gz9:�%�˚���iNaP���x���.����3&�r����6�E�<�ա��~�	�N�w�R�d|��̾��:���	BZ
�I3�E�9�F��H}��:��<��ER��g�_�l+^Z-Ȯ��V��
�w���NH�[1�'�ϴ�6�ޠΨ��8�?x��$}T�ʛV����e�}�ڲ�~���W���
0��v�a��\�E>�3Ռ|�ʞ|�x�3h���2�$`o�G�LT��O<G�)�����n>}_�W*+���i�ٖT\�^�2蒚����X�yKfQI$��P�����]n�PϴX{��'�":A�F��_���喲�+@���p���BV+��`��hTU�/d���(�yx]o��|��<��кe�ʎԌ}��<p_u�m�ރ�]Ϫ�d�	52.���u�KEMh{DTT����|o��rϲ~�vrd|�-��ͳ�/�ʱ��ӛ	#���7�$5!q��ț�	��������z�An@L8zF����J����h���D���tS�>�T��>��^����Zf�K���!��j����yY�K���D#�Q�O�b��E/6��R)��N�e�Bt}� wj�����E�!D32��"Mg�Ϧ�/�d9�D+�뗷ig;WW��x�}OF���}�T��ba���~�����q�AS�u�`�G��g�ҽ����
8��dh����cg�y筏wx�m�˙��x��G߄�ٽ��'xG͔RL+��w�C��|�>�6�Z��k��yk����UX�H�o� e���gg�<�t� O���'�t���~'>�s�_Ѵ�D���2`\�m��!�(��!=�g����m�sZ���i���b�v���g,4�;�����)R��ȴn/��_Ӱ�=#����{k'��������x~���/ի~���}9
���IV&�>�
�]Eʿu�P�K`�FO�������� /�Wޱ��"���ˋ��ksѕR etFޱ��=�����nΉ蕾��տ�v|�_�!��U&���s�I�����~Q���_>Oɹw�N���T�-��ߙ���{�Wmwp����!Q����ȑ�@���n
���G�����sЕ2�%p�*��n�<O/XyQZ]N��g�-�D%EV��7=�<���{d���jv�^��s>��}����꘲����}C�DwNT��$�jB�}����g�;	J��j��������7ܛ��nv�{��À�x~ɺ�\�_��>��nd�o�hE�����9�I�x8�,�+��}�����v���!��P�p�0;�g�G����]��ߗ�4T#���������qU��������z_�au������9}�x��l��jAϒy�9�E�0�M�.WB�w�TSD�c7�y����5�Bk��&-�Qs��B�-�W�j�޶��[���5V��Ig�9�r�o��;ΦC�(L��.�tq�|��LFJ�vR��9x������M���q�;?C���c$��Ì�#���z_���`�|~��Vq"��Vy$"�O[����1���^�i�tC��Wv�7����g�5�Vyl@�fuw���r{�gތ���{����+�������=#�����k���3{9�sC��VVo�_�%-�8&��z��p.��H>����x���ܷ4['�p�>0giDGW�%�i��}�~�
0�+�3��X��$_@#����l3mo�񿗱|A7��Q,��NyG��;tk&!������/��ޠ/�gVf���ݾ�QK�c;I H۱B�8q�����<���~�m}ʻ�Tϓ:�8������wמ������{�|�P#�>;~<�35��Y��\��4��1��vGųȌ��G<��)ڬ�LL��\�$�O�Gu\�xu:q*^�@Hxj:\���0q��p}{?������ˊ�4_�u/˻���6�0�h�H��n�Q�v�;��mq{u�B���X��m���c��/�G'9M�u۶ݽ�����©�5�ɳ!��AŨ�w�w��vB�����b�_\��{8]�b,v1<'kcӋnq��rm��9y���bիt��ڰ�yg�v1Ƈsn9Kq� h�g�=��E�A7������ŝ�0l�����6�/f���K��S�8�ƤL�s�7T]�;s>�|�����ߢ�.�oR�;Ims��Օ&�ċ�����:c-��ޟ)z��p\#�w3�Z��[���4��>U��y�q{��"����f�$�3�?[[b~�����y1����lZ�ϗ|ީ�&��={��w��z��� ��u���4�F�$!��֢>^�d}WB�T&��q����N�})�2Q��'��]񥻴��;��k�2=�xt�s��ju�`��ܾ�� ~���?ߎ���!�V�HF�����Ɉ�#�GX� �~z-��.o��	��{�v7��-ܘu���@ƾ�#�'�ｷv6Gl��A��?�Q1{���l���~�;��/��
"���co�C�-g�1��^X;/|;���D�{~�\l6��L��Wd`��l���49�Ի��&�J!7BռKM)�f��)`����j��v�?�^����f��~�flf�G����}��O��w�9�>m}H0��2 �����'���}?&�/�ۍ&Ә6��L�!���떾pn7�m��A-�ܽ[�F�[�&���7�9/E.�|���ō�ދ�UY��tg�*>�'g����1�D�=-1 `�{9���tO��D��8p����}�;��cL@���^�6���DB,����	i?	�O�Ϋ�]�o=g�)�F���h���GN2&��-�n!"����?v��4z�u����ML��w|~@��t�5�����m�#���a��!��2���ŨI6 Q�}�E }�;��Bȹ�o����p7����Y�0�"�h�Y�Nk>��u�D3`���1E6�J�Q����Q�[<Ɍ���F���E Z��m��˭qƲ��}� +r�H��;�>�gU��������~s����%^no&�.�۸����?AQ�����E��mJA!S4�:QU�ϸ�,�d� ����{����$�|<0���:��E�a��^1ޮ�nu��>��p����A:xC�q�Ȍ7���YJ�dFVbS2owri������1�k&��ݭ�kr��C1�e�Ĝ֣��c�HS���ۋj�S�����������S�ox�`���!De�GJ����eȖU닝�5��X��Ln�#$C��/�\{	��꬘�Jȁa\�e��x��_
��ǝ��Rlf���ݬ����g��U�f���ģ���Ї���KЃ1�-�_,kx�:ETAQj�h8���S�fz�!J����9i�K��ß_hj���j����r_N���a`�����A��ԏ��2���&��jǨ��>�>�y�k�y�cE�3����2�w>+��2��GTKKl!�;ˣ�]7v�/�dǖi+|������������h��۩պXVqۚ���2�<��.�x?��ʔ����xo����r!�
��]��Ճ��Cs��xm��U�b�V���]���8FM�;���
��K�������W_^���&�.9N���93�Z��g;�}J�׸/b�Ӝf��1�y����F��>Y�x�v� bgB���qX;K�o'�G�#n���tC�K�oB&'6��4LԮrf����8qf0Z8r��
{f����f���}f�}�OX�O���t�G�9�1k��%p}3�{��[_<�D��w�O�R4��	�:v�fc]�g��ݬl^~P���H���߇�˔�:�7���.gwO��[�>�;��HP��ճB�$2e@3��ݹy�b����색v#�\أ�В������Ș��	ܨ�޹�n���$u���ѧ���1�p(�|8[w�/��M�]G�QM����',�.��w�i]�.\�=��㭭�}Qh���m8�F��{��GUF��'ӻ��s/[�3�ɥUӹ�T"g��o�]֙�$��j.:SCk�.�`>���������9v�IO��ٻj#�{�p�c�"�fa�bLU��}Ѓޫ�tW��ǻ��qRt@,������/GP�O�=g����}�Q#o&ތ�!�U48�A��]���l����m��3�p��7����{�7�鬕�ZF)Su9M�]�za��B�m.�Z�Z|'�Wt�螪���o[8;#�U��ç���S�Z��7� �3�9`A���|DP!H��@��_}R���6b8G�"���5Q}w�o����1NJ>��!�A)x����d'aM��%����#��^_�ꇼT8b	(4`��do�����[k����z�~�!���K�p.|y1W�N�+5�u�L�/up@�#-�؈�z6��$I\�S������Z�i@�rsY�_�-z�v�T��D���k�~o�7� (�2�H��|Y)�K#f<�t�Xҏ]�&4�����(��bA�J9��^W�����b��2k��íOn/�lr����H<>��."��rx�?^��X`���N���aW|��[��r�$�Uu*����y��i�O�gĜ���R�ur?1�)X�8�n!����9��v��xk3g뜭k��9��TzF���QV�i)5XȘUsj�3����s'oU�un��<�Al��;�p+���t��{�G�*�gz�
���� ��A�D�}^�7����l�����	)��X�ױ�F	a�1 �p����������54n~Q�'�*����օ�;e�^Ͼ�v�)�SV'��zH8~>M��k]��i�3��ݻD����㐶!�*�`���ns{�\�����Κɞϳ��oy��#��97ᥖ�w���.��A�F���ߴ()i��-���7�+��|v}=5��e�m�s?#�#�mF���I �eL�%m�D�S#��B�J�Ƀx��"~�w������,���hN	9Q���hz>�b>�g�c=f#{����o*�1��߾m��=��w_cK��h*�A�ݡ�?\|�`������7�{�/Mǡ�Z�pT�Y#C����#,��w��!��c7���ځ�J�C�}��ϟ�F���";^[��O46pX!h��")E�=P��ܪb���(E�<s[=ϟD����	�Y�mΘ��t��
T�k��0^��fB�=����)�o8�u�5mg�W8nҋ�tĪ+u�8��fz�� �ݦۣe���;Y��5>N�'�\k��H�l�S�9λ!;���خ8���w]�4�^Ӫ�8v�χ^�.{���N{Vt�7���v���k��\�Ck�g��;����,u����R�n�6�|��n۶S�n��K�r�S��.��<][~6u|a�q��1��UA�N��g'K�������T���=�d��e玏5<ݺ�dst=�h�YV�4�~��[���$qT2���_N�	Hw�h������Yt,���f4�^0+:~�{A��bfJ�"�<o�Ǧ�����x~�9߉��ޮ�_y����W�_�s�^�K�Zڣ������1_d��_��Q�Q�a��'Զ�.,�����W�۞��� T�!eM4��o�}_�~���3�Ln��	2���/�z��1��Z>��+|��d:.lB��H���{�}tO�1�(t�~��f�`(�x^�}?d?���~����pS!��w�;�,���������NzRu1�̹�Gm�����d��v��ݠ|�����	"]}$�B��sY�.��z\pcL(�׋���6u��K�����߽ދЖ ���2q�z_.��#n�s�Jԗ�}��Oz�)+�gL�M��6U-�<)��΁�8eO7Bf;f�����J�%���² �
>z~K�UUD�؈�Ý�|>�}>�Q�����q;S}�m�t����C�7v �%nf6\WU=2O��Xh��Έ���X�"5Wu����>c���$�j[5��|S;������u�X��$���3k�_R�C��z���us��37���yv�`��'�}H0.��\�A��q�W;"pK�)5a/�R������#�H���"������>���_&�}H1؛��j-2�L��h�w-�ڱ�5��)+��źb��F6�l7RK��&.}�ဗ� ��܅bw���@������ǆ~Zb+B�!8F�Qq���;��C�~�z��i�m���)�e$���
�k�=7���D@;U����3�_	_V�'U�ۑh^���ҒF�e>���r�DYˠ�:�s�1�K�i���n�x2uM������*5����ySaꙃڮ���?5���}�N��7u߁Z�K�2AR��v8�iqx����qχ�~:7~���wS����Z2�[Ej2)���{7�rl��y� ^1��޲��_��=�T�D�ޘ%")GB�^���GG	�����-?���W�i��VưK���}�I�6b��O�&Ľ�����T�r�Lm9e.8D�Y[Qu�r<����w�&���n�D(��_-��*Ҹ$��V����o��J�������ook�OY��榐q{�~�|�|{�6�  �aD�+�4������[���y\|I�?�f�Ǩ�ߊ����c`�}�2�S �t0\(e6���o�sf?~�$�U�}1�:D?�d�T{�H+)a����_�߯ *	"���%i��N}�v�I�w��|A>����e��X�&,h�V:����3��c�w�il�l�n�&���)'IܷV2 C�KtVR�37���c����su�iptòjv�{��w�����w�۹�p�|j�1��tmYf���&���U��]e
�nYI*3��~�{=����v�*�x�"����Q�o�}�&~�,�{��b�)�AQ�F,�q���gh]׵�͗.��v{r\7ʹK�F	�)D�P�)A����*��n`��cd�;�HA�}Y�WٽCZ��y����{�y�w���V*X�OkK�}��C%f����=��g�����b+z���ЧN�+��E�v�'�l�b,2�<�"F��|`�]���	H��vLϗ|�(	vz�����t>�`���8��P.P-�c��O�zg��v���4Nw����{�¼lZ��b.G>�}\�wh �b�Go%�aL��Ap�+�(�n�A�����dp�r>��;7�tc(�'�f�Đ&0�������X:fElʉA�[�W�'���A��8; �c�ؒN5}F��Z���� �y-刨.<���>���_��߽��\m�u����y關����l�nű��n�FA�P��=�����ɱ S(�6�'ɭ�p��5�����w;�;�q�׊y��@48��X�xZy���Gk�R�b�>z�i�1ٶ��ϭ ���>[�m�-M���	ث[��ہ(q��g���dw]���T{��`�0�U�Ǔz���$���:I��u�1ф��\��v)e�@�A�ংy�k��/y=���vۦ���BaC$���h��달��s�v�1�ڲ�#
ݖ�)U!�3[��ڻ�p�C^63�~��S?p�w����O��-R����3n(�$��G�uf�
�QZO��7=�z��7�l�BE|&
G��z�b	H=�nw��~�u�O�4Ik*�A�U�X��p�/e@�D��G��e���{�/���+��%5;z�]څv���p��}%���Ly!X���#�֙$�h}�P���yWR�K�`�:ͣ�p�V�V�"~���럮K��;����F�������P0��=��o�}��\�=��k��]/����4�FYm�;�y�U�(�kv7V��p�DRc��Y��,�L%,�+3�������M^�OK�[ ۝��.���L�f�|iX@��QM��8VБ�"^]��������=[��D�C[��;������Cғc��_�w��q>O�W.���g[�����цէ-fLaZ�-��������"'{���%g�*�,�gD�Y�$`6�>���f|_�� �I�k���n-��Z�s�|��:5�>���,���A�>��/��z,-���!Cj�\q�A$��~��Ϫ�3���Y�J^� s��C�1����<���o:�5�!;�Wl��E���~�}K�|��E�&6�h%x��',�ȁ�j��};'Lp1BQ-�i��\��W7YR�<�<��ۛFq
ŧv��ݯ<G4�F���.����U:A������ ���t����௤��ln�ּ���i�i�k��6�R�pm�"\�_<����}�ގuR�B�Q����I1��"�q��K>fЧ�3_/F�i���Tu?���F���8p)$E{��>�*OKg��'*��a�?�=q#,�&�w�ԉ�W�<8���9G���<�?�w�_{>{*�#����~u�[�S�|~���C�ɐ��`��0`��.j:�P�>=�����"�+��'�H���I<
~�*�ʴ�����췣7�럺�x�Mǔ\���}�����鑵�זOy�m��4�:E������P�U9�igXN�A�8$�(q�!��DK�)/��O���h�!�g���:iݎ��Ev���v5�v����g����O{;�]�����{^��e�{��~B"��a藺Z�"����s�ޫ�5�����(�k@3�ܜǿ	Y�w4>�p��f��!T��^~4'�E-c��*}�+����7�QD چ��+g��cܦ}�2e� ��7E��w��V��$P@}_w��P��6�|߈�Z��m!\�葎��l�H���2F �j��d#[��Г�x��6��3\��"g�s�����]�|��n�@�o�z�,Ǉ�ts�pm�wI����|���Y�+�s2�`�_�$�8����H�w��R�#!i���_}������ܻ�l:c�%|G��n=տƊ����iu����?~�i�>���TE���=u��債�7��Ճ�5l�D�LE����r��Y%������쟴���
=��O�i|7Se�F9�P�y�vL�#��������+l �Ⱦ�s��7J�͇�9�0�=�p�n{=7�g�ȏ�k��7��&�VA2�NE(��`w��;F�	��P����ɗ����(@Y����4�M�*
��P�4�Q�	$W�V���ެ����Ǳ}︂�����J���~.��ߦj�xsه��؋�\bI�	�ޝq?sͮ�4�O5�D]�{S�]�Cs=�|I��G��g�)������|��6%o�C*gr��{8km�N����u犉�)�d���ޞ^ٸ
U����wk��ƹ���?�#�#�����N
��c��A_��n=s�aPU1�d2!�gQhA@@�drP��7�5�*�kX��B����"(kX ��X�*�*"������S�6�_���B�X!����ٟDq�a���P��>��w}��o���>��8M� 

������M�>c�@�����AYe�A�?��;���#�hX`�C�C�G��q�>O��� ���=���0���?:�=�{r?;�q�Ϗ����7yxwxC�N�{^����}1�+O	��?����z:������?���t>Gɝun�Yǲ���[x�4lL���D�l')�X��n��Y၉�HD��a�/h�m���gU6IN�Dy�Q2��p���D�4��V���m���#�:�����+��;ik�����H�]��3_w'�h��b͎�rě���k�-�OI{�!.�8���btX��X���q-��ޚ�;�4�Xr�׺�'�F�e�L^C,j)"]���ǌ�H��b��}$��4�ܿ�ǫ]����zC�MЦ>5 �x�z�  \��nu]n�!�ōbc�7���w�]zcY�ސU�DJ]�@��+KS�U�q;Om�9{�����`[�αu��vos�Z�ں7���Ŭ�7��"�u�`1;��kR�:lE�-��1r��R����®gdU�͸^ve{�إ�RPY�w/8��lzp�l��w�\��kmW=u�����8*
��, 4%1�"D�4�ߚ̸LAD-)$1+!L�HD2��Ҵ�@Ҵ��4�BC!1$�AM���C	HQD�PPD��E%%,0PҐ��CHSCCM��1K@DR�DMLCJ��$1M4�!4�MЅ1$�CE-!$�M!C���10C�211�3L�CLC��0CCBLL�M-	IE1�CMLCP�ER�%13344�$���L@D�4����M44���0�1!@�33L4���LM4�L������SL3L�LLM1�ICL�LL�0�14��0M2LLM���1L�ĄM0LL��S3L �đ,LLE�1%44�M10M1$C����C���14�L330L�$��2��14ĐL��3DL1HI��0M4��30LM30LLLCM2���̄��0CL���LL�132L�0�2���330L3C$����2L��CL��30�32L��LLM4��0LC	2�3$L���@LLL�L���40���LM4��ILL��@D�I$M0�-IL31�331$�33�3L������!1�0�314�3111���1332L�3�12LM4�3��L�0�0L�L�L�($�$̳��2L�3L�L���34���!$�0LL�3�42LLLM12�4��C3�0��$L�3�A1%DLD3M0�0�L�HD��4�ĄLHJ��M!C44!ҌH�,@2�0(�!JA 4#$ D S!00�"J� �2L�J�,!�³  !B�"� L1(Ā@�)@L4�0�J�	@4B� PP4$�J��2�H�*L4	@0�+�#2�C	0� P�
��"D�J4DA�B1	CADJ)*�1*L��JP�H0@�PLP@4-DP�4@�)г	JФ0�P-(@�ȓ"D"D)@�1 P�%+�pE0R��(h�`����Rb�&T�D��
@�"�(%B
�
$�&�(J&P�(Z��R�H�!J
V�a
@(Y�$�(����i
 P���������eH��ib((")	�J �h"��!
d���b �(Z�%h
���
P��	���Z&
�b��(J��b (��%��h
V��&(B����I��!�(��������%R((�`�P�I�hJ`(�h(�(�f(
iJ a��h����

!���e��H�(J iB���I�((��(i
(����
&P�h�&��h�R
)hH""� (�hZ(
V�(�h���R�����hfA�H(X� �&�`h�h(
"(
	 (��"���
(h(J")$H�������")�((���(�(&��("�"���&�)�(b�U���
������"�"������"R)��hJB!"!)��(h�(Z "�!h)i��
��$hh
��)j�`�)h�f��*j�j�*���Ae	 � ��� �h��j
B����$��Q���"�f�*��(�$JF ))
(��!I��bi�B ������������h
����)
�(B$R��h�(H�h)�R�P�`((Vd)`�ZF��Z���@�R$(�"P�)�)"JR�h��(ZJ�!hdF�)�!��@�$	�("�
�"i(BR�"T��Vd����&@%R�ahP��������R!IP�"@���
`����V �
�&F����dY)R� �� �(�Y�Q��I�(FE��
�D��B�)F ���)�J�e(��"U� (iF%X���(B�((`%)hH�)(�(��&�&Q�A�E�Va��	���	�
hVa���hf@%Y�X�d�`���b )� �hT��
R�h�hi�
@ ��f�D�	 �BQ� �@
���dV`@$	�X$Jhd��J�@(V�() �eZi%)�
E��i�@$��If�f�!
h�$�&
�a�� �hR$
XA��f���	�fT�T&	RT��H�d�&	� ����fY�&d��d�&B`���!�"�""�%&ffa��f`�fa�`�F`�&	�d��`��Y��bff`����Ba&	��&	�da�a	�fe��fH��b�&	�ff`�fi�f�f�fd�$�aPbH�%�I���"a�d�`&&	�d��	Re&Bfa�fbaf$�"B`&e�"X��ba�bX���a&H�� �be&`&$�H�!��	� &R%fB%"Vea�e&e&Fe& & �B`fFafB`fV!fRddf`&`I�e&`�a�a&	�&I�e�b&Hff��H�!��%&�d"bD���f���&���"X����R���������i4:~��1����_� 

�.������������~���a���:}i��!�����O�}o{�A\}�?�4�n����@��������0�ה>����P�����}����?��~~�^�>����_��� |=�|�~/����gO���y~�1On��ϵ�~8�h((+'� �����C�������@PW�z}�pc���i�v?Da���L;��v�3�t`��t2�����=�;���<��T����'�:x�	  ��ǰ��!�g�����}���&�O@`�#�P����_`����c�#�}Z^�����g�� (+>�Ї�O�}?�� q|�O�~�>�gg���ހ�P����g�I���C����~����^]��P�4hpg����p��#=���}π ��.:��N�㲞��Ge�o����^����������S�{�S�����&P6�����=��Ο�=><~��A_�}��_᳏��?����>��a�3!�c�7��Ї������)��Qk#�c���9(3���{��_���1-߾�   t                  
(   (     �      '��UR��	*�P
�@
(@QEPPJ����PQ@ Q**��P�UI �=��z��ʩ���Z��ɚ�5�4����mj���v�t9m��)��u[�lʥJ�4�XѤ��P�[I�p�"��Q@P� �� N��J^�n��w[1���ݫ�y�K�L�xou�J7wx�
��s���i���ۼ������=PW����qitv�wW��� �� Zy�@��ay�U��9��ׁEb{�\���Κ^��|���쐼�@c��Ǡ��׽c��h���C� ��3^&���I"���*P �@UP
�'��΀��;�C{7;��1�M���6mn6{{�n��ܽc��%-� E��R6y�<{�QR[��)��zo!��y��{b�'w�w�Tqz�))xƕp HT��*����ۖ��d���
�nS�R�����e[�{�D*���=R�:m�֩L�\ (�{jH.{���U���y4�]�y��Zҽ���!E�	JP���@@P( �/^�]� �w��!�xû�.�@�u��̯��;�p�u������^�=(sk�骧��z�0���E�\)x��W����gW��;�*�V�������w�-���cTNH@R��fM�I9���Ж����c@����9��G��ם��.��Y��݂&�n�ٵ�]���J{g�}����;�Eu��|�:��XQ�=={[��7��Ɗ*�t�@'�@��@*�QEQ%=��W 
����i��=f�5�w�����W��Ҕ��}��W�`� ��=I[kZ�s����y��bS�o,����4�0ꪪ��zٽ�QW��]�I�ѩy�����(�ѻ��︾���s�Һ���� ��K��G�"w�ǭ
��â�{ܠ^��T�ֹ�{2�p9{wc}�W�����Ž��p�B��*QD�ptw
�ty��E9j]/n���w�M�����"�z��!=n��/{GsR�9��=��v9������N�v;���� s���=9���]�=�U ��4��=����4�s��a��99�As���y��g�z�H9�pP{�TQӼ����W��r�r�/�  P                             �(j���SJi�'��CL���b&�~JJ�       ��R�OIS@      ��R	��C 	�   &# A'��L� Ți=M���4ڌ Ɍ���A!��#4z�@�  ��_�����k���������W��%���v�o�ն���ݖ�+\�������mV�۔ڕ�}���[[V�w_֛Ww��;�_ם����OK����gk����o������ǹ����n[��|�����{Zڶ��z��P�|�kj�n}x���-�o���5��҅��t��_�	 I/�b������կش�~�����[! I/኿���K�����E�4HI/�������l����ɽ�E<��͘c�g�b�\�/�}`o�!�r����*^{�x9ݶږ`�C������&l R"Cu�5T�9�P#^��ɩt���ǄIh�º���oe��6]�3'����&ȱ3�D�-�~�>hₛvof9��tY��9�J�=4U��p�oya�
y����䓺�sjX��d�N�v`�p�G;�f�s��]�^�G-�^<��*�{�)��Y��j��Y.��]�#q��ݷzf��ҙ��'vMA�`'���^�t5m���O.��f��<���Fx{�x����[�8{aU˺�3��:�]2]���Ưwp�3y�q��ᜃɄ۲w\RɸpC����4iR��\g.�y�5&r��q5^#�wxs(G��U�{H�B�*#5ΜK�ё���w�DrAc9����w-����i����UB��+V�W���f�b���-tK�� �2`�!ås�Lx��6@o��n3�������5Me%�c��:��A�G	�h��J���ȼՒ���/�BR�t`�sN|�0�UB>������˹e-n�x�܇g׷ꮰ�x1�3���ӏn*�у{�]y�X0څSK$��6
��.�a1�zZ��ڃ{ϡnk�ےjx2o�G.أ��OKW�2�qc6���N�a}غfW�C\N鶾��*/v����.�m�Ӻ1]�y7J�-]]3KsJ���\����T���g���o}`�ۏ�b�g�i��>r��
�ӻٓ��Q8hS��y\渳��my�L� Y���� ��k��G��[ќ�A��x��y.k�Fb�Ș7�#�Uot���]-�ik�כ�Dg�k��ü7��ܖ�׵C���׆�D-����%�c��"�J%]���1����Q��,]���zy��Ǚ�V�Ӕob7NǑ�\�U����;�K�H�s����Z��˯;O\�5�\N:�x��8������.z!C[�����׎���˚�m��zV�����\=��d�3��5�kV��1ћ��r\�:7,S���ؖ'Rd�\�v�Aݘ�=�e���;WI��Gk��5�.���4�u���݊;L��ukňd��9��Q��܃h8	��w��J#������%����SA<3� ���s|���9���ӧw�A�Qf�������d��7w{�wb�iOqU�tˈI�D�ǃ)c�+:���B��u�����`�D��0���P�f#�}�yb�#yΌ���c� ��'lk]X&|�Ql@ރ�ޙ56�*9��8��M�r�{��YGPVjÆjT����`�3w���ݿq�zc�v��%�D��w=3�n�{K�%">��6^�uq���_�u�^ņ �>�,��9�۶� �ܭ�Іa���?�^��3�nY0��^n[�Vڻ��`�Ij��5�u(�i�u2Af�u��Ү�9��(9��,Z~�����R|jݢ*�,���ЯL�-Ss9�؛*κ���:�)�lͱ�*�\�������4^�xI˽#֕�Hf��r�:���{7je�wh�7-�C�˗EAv�[�M�f5�c���xD43�%;u�m2�)�W>79���[1���볥+xr&a}S�h�s%��-�DZZ���t4��ݻI��qƬ6�Ǝ�}ݙ��9b;ˈ�մ��m"t׹�gktR�48r^�֚�A�X9��x�i��=*A�6Y�G W��]��$	#�`�rY7y4�Ze]�e��Xٔ� ��C��q�ۥ�gL3�iAZzs[vĶe��cX�
�y>�����P������Y�z�7�^��u&A��w.�Y6��ٽ�ý9�Hy��"z���<�4�c�D�Z��+�Q̻.&�:��^I�m�v|y�Ի\�������7}mYJ�3��f��:]FX�ϯ��V<���fo�F8P.qG]�nj��W�b$�M���d�9>�%�`��#pj�ugoQ7%y^�ׅb����Uf��M\jY�>C�,]��0EΨ�&%�4�\9,|��8%kse���{Z�f�}��ޯx�l9PW�h����X0.�m�ݤ�~���ŵ=��tɖf�ܵ�$����"�.ㇽ�ϔ���ݶ��ՙv3.{~�Z	��P����#G/�wc���D.����+��x��1�5����w(e��]�[���q�n�	>�Oc��C�����.�êe�s䳲gaSF
99gt��'c�Or����cŶ�M9�6J�g��k��B��ToQ�:qP��ˉA*�J�X!�v����w�ɳ��h��u�t�N��ΙۃJa�5�G�]U�^[Y�v�N�v�&��(U���_S����u�M�9�f�8l�{Q��xT����˽��(��y,��7�{�݌XG����oV��'B�c͍�#{>�������Ī�f�z4
�8��
�f20J��q�U�\��c�r�3ykp�s>��fm7F6]�&Eh<��]8/T&[���n�.Ӛ켖����o;9q�+{�g@W#݉���;�z��=Db��la͊�	L��lʛX^;�5g����w�L�Q���{׾1��sǚC��{�0�|Y� �7h(�Y�c-ܓp˜�"�fC)�uP��
�+����V���Lc���3�Vj�c'�ɹ�7���:6
��+��s�ף,�6���ݳ��qsᶤ�Z��b@ܻ�N��w�wF;N��l�wU�L��;��Ҵ����tbn uj�O�ٷ�������<;�+����6lo7�������-̷�/7��,�v���L�����T{aycK���7n�wH�wkoh�[��Fo<�7��\�,��A�/y|�f.2Y2:�l�&H���=ǟv�(�Zp�:����d���,/f0�4��<s�<�<�^U3�LrG�k#�;���_�B¶.��bv�0���t��@���q>ق�ۚԛ��n���`/�7�yf0��Ώqv#7v!�שg��웻�W0t73p9ٔ��K�#���"��&\�F�5�����z��va౾�%��s����et����'�ܞ1^�{ob]�8��݇�P�2��L�g�y�nwu���n�����8��O�ۅ��F`�u7Ӧ�L��۩D�qh�z��B��nd<j�6���l-��U"�#y�5�B��%�W����3�x��u&���ȉ�nX2����;��yѐ����a���B#O>���S��ե��H�nOy����I׫�ec7O���sK��-}���~p�7M�ޚ&Y7%;�RuTY���6���:K��^�;\�WN�F7������]�/K)ˏJ����݌�hǺD�ϱY{��Q����D�P�q����oJT��Nv���o�ݓ���^��,�Òǎ����;H�Yr
��Hbi95��p��I�YP��]�D}{4�t�w�=5bAK|���(���eőﳫ;�^��(yL��J2
fB��Xq�t��w2�����+277c^~��e\�6�Ƿ����{^�U̻f-q'&��R��&�m�$��ri���^�b�r-�;��gv���\,v"+�`����ٝ9�ݧd�N%�-�R=(aS)iw1�A�LS�LB|��bY�,\0\�sq��v�4��v���0�#�����k:�&N�*��LD�����1��gj�nq2��&�Nr<���3տҼ��H}#��x`��d�x����Fe���0��[���c{�X��z,���tsKx�cI]�%��y�U�b�v�NaR��pK��� �a-�Ci椪;r(�7��>�\b�JQ�|�eڸՊ�Z�<�}�z��7��,>��H�H�a9�p��["{��2\��[�������0x,⻸����}�Yޞ��yZr8:J����}՟+ϻU��\�S���V�;ۃ^��`*��f��
�`����C	�h�=;�ǈ��9�	]���V}�2FF:�w}�F�ݛB�n�����y!(��F��&@�ܶ��u�����?�fO^����Q���v�WK��=�ۨW�;wNH���3���e}nn��d�]�Ek��n�@��'���ư�Rv���8��������O��y�?B�yf9Y��z��7��}�O�{����R�
���S7�y���ʛ�W��҈g��v{<nX��Z#�x{n��XV][��{�o?{�2�
o�A�)u����	HƩ��coꋏ}��:�bv��D\ ����<H�"���;\;=�5!��z�mѬ2��y�����I��v��oҮ��'��ٞ�{2b>��z!��/�n�;�4��dkj����B���v���ļ-\�|O���2`y�'���E �[Q����P�f�<�)D���,����q��yv�/)���^f���[�8��SJ�o��{=L���E�ۣ8A�|����oJ,~<#;m�Xr�m�]������ewsbR���<O�U��x�'��w:Sn�L��I��;�ķ=廝��e��b˻�곰��섞�nt��򙫏{<��y>�r{3c�olWN̽�H�d��<y�;�Td}�f�xwlb]�N骫���������~/�F�XI^R���E���UAH&Y��Y6(ۿG�6�jUH��c�u��T�fd�~����yӚ�M��.l��z������s޳�^�n�3�hr�9s�Y���K+���a�QIvf�{x�f��^�t퉽ց�j����Y�F��O7!w;�a7��;�����+���M���Q��%D�qM~����+���y��t��{v��%�o��J;=v�I=���ms[]*�fa�-�d�ɳ�G��J��sF�_g�Z�{H��F;����شg����x�;8PFa_3���*���4]kxNz3r8*TD₆��Y%�R^l�V�קq����$�s���;�q¹R-�E��~C�O+�]�;��m�����9�)��_(�3y��%���Nb�+�L�/zݢ'���)�)�{�Ժ���L�X�v�nNy�t����lsR!�U������0��wVOON�.F;�l>x{׷��.l�/��8{za)���a��o=Ι�E�b�4�h�U^n��<��<:z��Yۘ#��]/z�3!s�5�v#��`�Y&hO7f�z5U�+lk�g�����I��g3f�Bn��l�Rt�
�w;n��5�QîdD�͝���b�vWVM1m����sVY�9�d�O���c�;ibd��q	�hn��ɺ-]���7x=��R�.��.]�zh5����[�o�,���5̾�9�U����sqҞ��D�fL; Y�;�5���7F�mȗ�oS�{���:���m�{�7�x_z2�E�OaP��R��o,�)�ކSA�i5I�:C}�C«"�uԷB�A�C�B���K3�hgh�x�9�-�	8�
���P�Z�DjE�8�����Z.���#V����Ⱥ�;�Dc7�X�電œ�tZ�K�� ���Q���̡2�ʒ�1������H�3k��)�%e�ɭw��-�sv����ZT���K�[:h�橈̻0H̓�I�r�uf�<G����8�&�����`Xfכ��i�u��qq^�;!���Ђ^+^==�}��''�]t}V	�f,1�F݋��q{��Z�:
������oNQ:��r>��W�"�,ӗ�8j!����m���/c�{^���E�}�8��ݝ�$��6"N̻�7`�b���Gc��W#J����#ٗ��=��(u�w��Aэ�L��дK�L���^�	���H���+����2�G"�9����Ѳ>4��v�.\3�eioC���/d�Ƥ<P�\Ǩ��ucW�4'Bۼ�;��:d(�=��B�G����c;	Z�����운�L����EKZNC�tŎ�K��Qz�ͤ�V��;�z%׆�^�r��G#6�Ԗ2����q�3r>�}�Z]e;��Y��Fv��xNy{��*���:y`�kU���)!M8q�f�.-/L�Ӵ��l��3k���vakC}Tn�ےoޜ��#��33`�t��2@�n9Q�� sB�'Pv�wre�vG��谻�u���"��A�2of���ܓY7zՙU&�rN��wf�-��f��M��՘����f4-2�
;�Ʉκ�k����J�|(ӻO>�v���#�ۺc.��;������6Ç�h�R��]^�6�p������e��E�S˧�o��.��'lU[c�Z/t�4�ke�b�˗ݯ4D`Vdo!�MBs&X[�S��	35���@~��������I�a��b�-�Y�!Ǧ��\Yi�RSսڷNZ���M���(��������6]<mŻܤv��K<w�3�<�����*ާ
�u�-:t�2�{s��s#�]�k%���s[��f���c7Ä:�r��bz�Q	����j�Y���ۿ\9Ǐn��9���Q�&[%�O�2|u��;(��hM�xfj�V�tì�{w0^�
�� ˪;
��n��^MO"��Z����Y��S���_f,J���]W�"��3PW�r`�|4fd�,��i��Jl�[�dHO�S!�%�R2=s������M9N2;=p[,��dwu�е��w�'8z}�=n�0U���N�u����M�r����L�7s���Wu�Qk��r]�p�/�v��K�ո���eParٰ�@��^%�R�/Ҭ��y���޹5ͻٙٽMo��h�����ڈ���*n,GXR�~)�7�y5Ѝ��Ջ��ɹVvB��>���2-y�Pfw4e��=�2���˝�-�׎q�E�OgcHfwh��ȶ<ۅ����˂�s�(���ő�4k�9f�0��v7��vNB�u;�9M�#p��~o��~<��y~o������H�%�}�X���G;�~y�M�N0��L%�<?���ﻏ�ٞlT�뫜�/$����t%#��
����H���M�a������2[jL�Cl� ��\e��lw�?�-��c��B�E\)�mԑ��&H8� L���cvy����6�\�}��z���C����q�gu��Lu/�gqw4^�1F�􊛇���q�����8v�]�d�]����p�m��A�U/���ߧ[��:�O,l���N}|v��l5�����q�gf�
�ak��QpG#zK�B�7q�Şָ����jg$�kZ�Ҭgl	IDh��d��:=�0�n�ط�b6�Ĭ�e���nЬ ��F���`���hU) �GVI�(ٚ��J�&)�j2���dD�df�RR��Xd8�i�ubAo����fٗ���k�Cke�ٷa5&N۞ �i��=�_u�í�#v�m�PsE��v��J�e�C���Ͷ6��V @kά�׭�����c�6���������d�7cg���串U^�ۋ�m��\6�ԭҽ����^��:�5�OKQ�<e�lr��;\Kn]y���q�H�X�<��g��N~������9�@<	��q/Yg�UՓYh�Y�Q���R-x�V�Q��u��V����SE�j�Nn����:�j�A�C�ᛧSvx"��`�j5��ui����ҝ/:\&y�x�{�=��l�j�ۮ^��`t�X�!>���v8ݞ:����j�v��ݶ�r4rv^�NՇa��g���.�A�,Z0É��Jq�;�v��]�ú��{y\ݍ��rĝ�����.��2�WD{�y���%ak�7A��e^Юo3ǅ�Y�2����t�{\�0d�M��eqt�Gλ��rJ��\���x�{F���g��<�H��9��L��s]��${6V�")̹x������d\��=�[�f\��ѷ���&��v�8�u얍�":S��ۖ^ٺ&�q��t۰&�j����gnck���I�{ �quȍ�\Avޱ5�ZT���5�K^��W6Vxس,���N�v����zۑ1�L��GQ��&�;G�ҹ��ٺ�\����)q���bG��GYR��� ���GVn�[��slܻu�9n�k���������B�8���pGQ�m��'���b��F���I���W6�)��.�)apq�ܭ��2��u�5�1h��;p&����8�5hl��:X�Zx�{cEқn8H�J�N8�k|Ol����6@��5<�3�R��k�{8����5�iZ�˛
pg�ۛ&z�����Y4LQ����J<���tqnc��c�VU �mAu�t���݆:��C��v��	�7:�����{&85���r����lOs�Ct�'d��hl��s<n����mzz��<����m���:��=���Ӥ�{l�{���;! �zs�f�=�/"@񻛆�
c��<z�]]�c��K8��O��L�n�glk,��[����Kpf�5�n��Ƚ�[�7��m9�2J]jG�"Y�V\�7/��|���;vx��STn@�踎�)�r�67O+�kQ���Y�=��{�"^i^+t0$P-[`dd�tv�F؝�R���;�f�{��Kt�뉺q��t��t)fm�kn��ѹ	�)����h���.Ju�<�u �q�/���g���v��r�j�[��;���Q�k;Qs]	 ����V,v�����j���78�D<N�������湜�ɻe��O+��]q��m���{p3��7 ������m)�T�+s̅������md�J!m��9��l6�<o:�쑮�:��ޞ�����v�u��f͜Ɍb��!%�(��zܷnum+◝��p sn���������)�A���v3�ms��q\���^8	{@'�� �,g�dFl�n[\���:wI��{�bF�k=�Wu��7X���h���{fv���ú��i�7k9�H��r�F�c|(�F҄��ВI��9�2<Oi�(G�u�,�F������ѲG뎁眼6�ps�������ͺ���da��Ǝ����M:[�R�cz�yKnŮ�]��U�WZEΚu����XϦ�4n;t����� ֻ33�cb��nܘ��l �;X������D4c��]gof����M>ku�����n�`�E��W]h�Z��!Tn�����(]NT���룟O(u�ϝ��{@�f(���6��l� ם�DX�6�WRk�����u���ی��@�l�P�7m�^᷃�5���o��5�MuؗkT�i�����-M�.�m��훆�e����tD�d��c�P�nۣ�M�on#�> �v�;v�Xlj�[�������G�h���qٞ
�uͪ��D�K+�f��v�a��W+6q9�A��"gr�k���v�Tî������|�������5{�,�3Qz2H�Z[��`�D��`����&1�n��]����gR��ܻw8A��v�԰�Ki�Y�Nyt�]��������7gn�n;��5SǞ�f'Lk&���И�ĵ�0���a���n`D�����f6U�'"�s���fy���ް��^�Wd6ݣ��f7q��,pܠ��m��wm�k�b�k�nK�nn��q�]q�.�7OZ ���\��8�ĪԤڒ�K25�Z�2�s{nχ��n�1M�=�\��CӰŹ��מk� L[d�k��;�gq]�iL.cx�y�洇��m��v9�Ă����m��ō�mUi7p�bgv�1�D�B�����}���Ԭ¾K��ƴOWmF�\��k.���O��֜v����e��l���^x�"���Ɋ�6�4e-M\sq���c35ir�Ԫ&	h�)tz��\�������atW]͐�]��l�j�}f�v��Vw�vHAZY)�ft��%3�$�z��N��>�94`����v�dd$z��`LX�i��lc4��Þ��Zx�x�Xw͇�6��Nw%���'h��e0�k��,�ڹ�,�z�V&
hkY��IR����4͌j�5��I�݂����v��:�ڡ�CذX6�w���j$��!�u��k�Z�j�<yJ�q��T��n�[�s�l\����7%��k�b�z�Չ��v�#�eV񽈹��M�v1�6F�<Aʝ��M��WnS�5k�!�g�Qܶ�;<����	E)][��T�U6qr�n�)яn0V�}�r{;d�;�ֹ�*�b����E�҂d<Z(h�8-�I�rݡ9����x{h@R�l��G[�n������Wve̗���k[��JWik�袸��n�5��3d�-۱(� d�rӝrulSV�����]Y�:D�"���c�ш̗ϊ����v�-��9s���p��#��wmuŶ|5l��7b#��2���U��$�[t)pe�V[;�:��'�I�I0`��v�.�Lp��m��f�8^�����k�+�&�+Lv�]�m���Wng�X.X69���W��4 ��xԺ]�=��.l>��N+���3��c��1&�bH\�bSl�F�u�k��A�����t�L� �[#���)�N�\�[�r68����H�@wgf�Gh�a��i�ܭ'dsv�Ƚ�L2Ն�k4 �[FsKvĜL�˪�v�zy�8��0/ew4��kQ��G�g�]���z�4v��ƭb���,F�
��vy3a��''.7F�c�	�%��Y�����ј'5�vL�s���Яi��Q�����j�1�rtޤOWS�	�FF�]:̰��:���ǒ׍�N롤�w�;�ֻK�vu�ݹ�� ���p6�x�=�+tr����b�+��<��q���KqF4�x�v��d����;[���Y�ɰ�p�۝W`�y�.�p�q�\R�<��\����2���{O���@�<��ڃ���j���u)׋j$�A��6	u��kgWFH��1�냈ܼv8�t�$�u�z�� �W���cM��]�k<�4�#�g�4ش�1d3�Y��$3u�5�63E��Hlo^�]��pڟR`��z0�sXfkZ�h�f��M���,�q��3��9C��[�#�&�:�&�u�W/y�խ�^�����s�&�D�:�fd`9�H2u]�E�_�Aў̅�3:w�c1�F�R7m�]���ZD�����u�w'3֍�	�}nn�v�M�3@��ubq�ּ;0&�nf�=�g��3�T�;Cbuo@Y�d5GE��붮ri���J�F�f�ʢ����]�������Sv�ژtE�� ��M�Y#��)s�h��c��z�i����by]כ�{y�V���q���捻69�l&�R��=��g���\Rdd��v궻�̻�W�5�パI��V�0Evๆ������h���9��u�u��Ӟ�b�Hc*H�1,XZ�Q��̸��n=��M���&��ق:�e��9�����6F)�8��H#l�n����K�a�h'�I��۩-V����h��]�FxT.У) �z�z7g��6���/�fd�d�T���SYڎ�g����L�u�s�I�8��3Ŏَ�[��%1�cm�X���`�x��q�n�h�&���C�V�	�+]X�<�#���V�q��pg&���h��[�|�me|]�=����Ǒb��F�3���ڎ9���Ʈ��W/��*��	�m�v�����&r��sP�aG:���+A���]��Y��E�K�����m�U����T�*��n��'�^[�z�pxj���'�k�M��"R*Mc�f,fn�m4L1��1�N�0�T��Q���<���,������vJ7[tnD1:�֗*�W5:B	6I��.�[�6�n�4% ���3v�K,Çvr�'�\��v���s*�^�h��L�!w7h\���e�6y�tƹ�K�oZ�Zm��d�Ach�F�fx#�݄����=�r����4fCK��]�ILGI�� �e�u[s��y�O]&�o�ѣ�'��A�v�h��d���}��,{D�m�Zt�6��`<�wh��3��r���f*:����ф���eְd&D��Lƴca��[�]R�ǭ^�W�BI�r\��~�����V�u�����V�oOk�������־z�w?�����_��}>צޟ.�/kr����Jh$	)Q���6�L����[�Z��%�%�I�([(�R0�d�
��_�`΋1�ܳ�H�	+k���	��|BH��p��>#�������)H�+v䦩�JJ��G�JS"��<;9ۭ�Ks�
��;o3c��[��b)4���D��n��S��������&�\��p4'�A'O)%&�`�}� Թ��)�wɛ��9��2%#.�=�sS�{��� ��8�z���};�# n��}�v����f�%E6�8�I{�KC�!��u/�pQWB2�J����5�1�u�#�&���z����Yq%�I�7!p��JIJq%��6w|�R������j�!�-F��y,KM��I8�EMĂ�)�)H�UU�������SM�u�����`>�Ɖ`�z#���c]��-�L����1q��3o|V��9a�O�#����}�z�xQy�(�����'��h\�.��z��ŏ8t�x'�Sspnց}.�t�����`��!�
h�(HlI���ē�� .�e�C.䎩����gs���ׂV �>�C�i�W�a�Ml�����ަ�N��8��6�P�eS��)���4s�ӑ����{�C�vwii�§q�TX^��������#(��������%ں� ��T1J�C�݊�Br��F@#OPD�����Cx���.�i�I�A�_<�L0����/����;D9���=�/�:���!�2|-���n��eTथJ�t�\/��v�^vbSJ�x�g�'�1�a��X(�� ���q{w�^A��75i>�>�p�ay0cEJm��UVEij��2�-�ӡ���7�oy�T��C��"�::Xr+]��ρe�1��{�a�v�3����}����x�OT��p��:�|�*��`wJ�-)E9>��h��2@���$�2�_;[�B�n'W��B���}ya]�xv�:Vߖ��0��|_�$��w���D�F����=n|��AuL���,���n겕X�QBorǏ�zq3*RyNn�&����� ����0��r���NP�!�z.�u`�Z�V�`���R��q�g�7S��X�7����t���;z�"�
����ŵDR�>_�FU<�ʽ0ʔB�G�hy�T�7g^"ECiӚ�������U�pm�>��o�p �A�����N�~�N�Op��czC��'�xv�#����wU��'>!e3��������^7r_����������K}}Mo�_47m�����J��(0�[-ؐ�Iަ)���u�����"�D	>)�d(V򴩾�>é�ȟ)ewU�r��i�Lޝ���4��{��J�媔9�'r��5#�?"v�#տbYj��|�OiJO�]�H�>��{|٥pF75�i���P�Q�z��pz��Dҧ���*�r��Ν�<{}޽w�ts�i�m��Z����H����V-'[#S��E��[NjMr��.���No��mi�T�&�3�����������������'!�o�Q\�"��h�
$�ÈCA�Z��{�)H&~`��<l*n��wKš	F'�Q��y�����3Z뽘��)����lclp��g�T�ɮ���%z%�o<��|�$��VU�w7�oA
8C(�+�U�]OHx�\u�w�G���H�Q2��T��7I�ܧzy���Y*�4H�|O<����7��g��B���Ht�V��<C8$ƞ_��Ȿ��QFp�x�� Aߥ�/b)h�P��+"Pc�gD6�Π[yx��ϲ��M~z��Gow$�n.����)Y IHtC��w��A?ae�o��2GɎՍc�[e�*4P5Z��	'TÞ�ۑ/N���x��#|Z?Iw���;��^�$"�sɪ�ٳw,^�����sF���Z�y��Ovs�^��o�K���&K��T]u�0'5Cu̧��;�gp�Po�W��_���cC:�)M��FwͩF��"�#�䁓�t�]<��q����J�`�g�xM��e�v������?"H@�S!��QW����
�äD" D�R`o�kΜ|������S�[���oS^��ʨ�!��X_'W�_1M�"!�����y嘮�}I4��@�� ~e�x�Y��&��$�,9��hy}u��ٶwwA�u�=����i�{�����.�M=y�^��#m�t&fe*�}�o���ڤ���J���p�j`e�䜩c^���9Z�B|�S�x���27�����%v&�]j�Ɔ�Nө���F��X5�H�9� 
@y��Jcf w�h:��qn��:)'�����j�0��5�K�����u�H����Zu�(�.t��97�M�ͦ��x�|��E=y��i�\������P ���K����W1�fi𦺂n����F;�wIHȞ1�(�<ݸK�z�.:Q��MF@!J�X�H6�U��6�-P ������&ެ"�dG{��	n�83�����^���+��uI=��:*�/���������y��#���W���{�d��g�Jm]<���W��jA��]��fT��&n�Rԣol'�1^N���E�0�C��<��k`������ԯ����K��8zIt���=�3���X��Y
K���������L�Ag���1\ķ���{�;��T�/r��d��C��zk�*}�M�^����ٹ�pʦr�wʖ��d9|��=6út�@���$93�?&��_�!'Q>?�C}���P�{�g���A�:=�p}�V����+{��j���71^���"L��P�wF���[}���r_+5�SЦ5w1�1*)�v�&u��xՖ�zn$jS���ĉ�G�"�������f�{����=�ev�c*���tn��Bj8�".;ݡD�hX��D�	3	IB��ܖ���@�o|���ȥq�廉ٜ�9/v�/><x���E5i42�q�Y�=�]��R BH,8�J#��e��<�\=�
s^�N�*^�{ַTb���X:sY�w���0��'�M��X�v�j�ة�fZR�Bsd�wr�O�y������JYK��2�+�����w���9�܁@�8*���b2�ʂք��!�c������`Êl�C�����p�sv���51�H۱n���a��� �}=(j���@bPt[���Ζ6�����B�I$�犜���#{�u׊D�o�0��K�EO���}s����c�����xt������vx��r�'M�����ǐ���s}&�����g�T����x��qѭL�8���3�2z���os,7X�:)5*�����*͛;�ʣ�b�^�z<?v$8�N2���̪�mZ��ݻt���v�+V2�j|��^�ՎG��x��$�	J�o|��w�(=�����2#��Ѝ�:��R�	AR����q��3Bs���9I܄)N�wJ����R7��]�J$αk��kz̽^�u�;��"#mA;{v���ZD�9�
c�^4+׹�'�00��W��{>��z�S�� pE�>�B�$���mФk�*Ҋ����IhL���kW{|�^�ER��W���{����xD�֙�ꪳ��'�^�>z�D�w���r^��MS墱Ԋ������`��$U�������N�/�*����:��/v9�]Q��û�������"���M�wF�����G�;�gyq��}�e=V�ܝ�4�Sl��Mj�����)���,׎�^���h���)cֻw��z}9=^����)�AOrRKS��
j��&J�Dה�s�p�])�z[�.�kn��]M���i��ni�bCh\ˮ��ƀ_t�q��~B�=gwb���׼۸]�v\E��%o7��}�w7�gNIѷ��$�վ�����bt�N:IQt� u�ĉ�T%uW�����w�*���W7����>���Qu;�Fq�gYv�ęmA-CWi)oN�ZCa	L��*�k��i��de`��R��3����:#5��D��7W�t!�Q�PD�Xw].���|�Α�3|��$t��h!lqY�r7���C$orm5���k���T�r�������U�>_b�e,j�Ew-T���=	���y���X�Q���<�%�gl�Ⱦ|vq�C�/�`��D#*�~�I�4�B@c�G��4	�N�!�w��O������"���f8�ʒ)#g"�"ni��a,L�D��^h9J��I�&�%�
4$�C��D� �&�Κ��fn����?B�Ï��V�H|�K/�|��_bx�ޯ*{H"ב"�u^�c"�}��|�����ᤐ��	���A��É�.�& ����JX��<Ԋ>C)�l��]o��"����|��*V�
0�����z�G�G�X,�*�B,$�U*S}�>�׹��Ş�b��_]�,�A�HC?8P��P%T����!�A��.�	$��ԧn&��TکG���x�ll�Z�'����yFVգ����)K������HaD�p�$�Pg��H��"����x��77����#=Y¢��Z5�U�`��]��������:k�Z�%R�'�4�א[������fU�\b����2�3Ȝ�8_aê��X�np'��y�t��o�N}W�Nw�w�q�$g=R'o޹|0�/3!������b��A�f!E��v���'��&J���V�֎�����ɏE�
����?C��7�a�q��vkq������FS��N��/Z0��đ"������'o[{�f�6����m�c�*L�������-�/)������,k����im�[���ot��f�x���}�؁�@҃HEb.;B��Ե�4@�BD%
E��0M���>~3���c]���t�/�,+�|<��v������-3l��ےԶ���2_^�a��6j��L܅��I).����Ԩ�/��F1$$	$�� �$�)!$��8�';�3�~��Lٚ�Su���6e���BT�7�δ;:��]�g�wn�vcR���t�E��Ϫ��lq�A����M(ݏi�6J7��x�.(ݺ��'�lz��u�N�cVN�nr�H��v��ܤ������q�"޹狂�ڋ<�G���B�I6�c��m��ҷD��;)������ەzKl�����tDt�o;��V��A��f��c�<\��c*a,\��G1=]e�lu�}�5v���.\v����x��#�д����5;����b��2�D҈E�V,�a�=��Mǒ1��l6�h�=�D<h��p^v�����x\Z��
��u��>t&��ۨ�r����$��/$q\]��Y.eRהc�!�Yn�<�؞,���1e[��
����4�i�m"��X�gTr�b�r.��1;g��]�ͯ�����A��V�:��R���#i�6��Ęz�m,�c��4�	l���s%6�E[Kw&�c��v�b�󚎒����<��a��N�=l7�zU܇&^���;�ܡ�y����m�{�AC�E�H;u��^(�1����Il�=�������8�M�d{�zz.{qs��c����� �v�L�$��,�%�!jV��&�)���=Z����.S����x����u��	�s�c��vW9G��lgU9��s�]����a�:�S#8ݖM��ɥ^�휲-#���&Ӏ���:kbS���ӽ�m9��6��5�은���v�x�gc����ޝ��p=�=����@���dzN��y5�Ȗh|d��ۭ�v.�M��u݌���"u.���Sm��Zmg���N2����IO����m��ٶ����4;Cu�ńGvK>�u�=�3�:���+Ʀ�۫�n9�l��n�u�n�{x�[���獣d58�aIpgv�:�{�� rf�6wg����-溷����]��p��-�5�^7C�����i�K3�"X�)]R�].K#5�9�t�pmb����y�]sz��K±�����u�	.ް&�Y�V�jNJ[
+��ɷkfM�śЕ������-���$�~��@�A�� gw�žOo;�幷����>� ���t		�$s�@�����yn�y/o���������%�D���9�ALzެIv��� U؄��w2����%�;t �UR��Z��l���k����֬@zD�� F0B��4$- �5��L����G���L*������B��Z��j K/(�q��{�� U�դ%�V9;{m��ު��Τ��J��BK��I@�c���*��B9�̾h H�~�B5�$����!+�k^��@@q):�:�F�&PB�%Hf�.�öan~�Dr��>�����z&�v���ܖ�7)	!R�:�v�<�Ù��#���g[^܈jx99����l k�F�UC�d���W�mkF������O9�6s�88�yy�aŮόm��]��sVO�z7��.���.�:�����r�+�n�v�y\hŨ97n;l��φ��&iv�cA�+r�JS6��d�K]gK׈�1JJ�7����_~c���m�{V����_I	ZL�"�a�)�	���;>D�>yTl�%H�X�ʤ��,�[KA�xY�Ǩ�d5�d�}u�Q���;B#y��v� �� ��T bf��f�%�crH�쓽�!�������n�rH!�m��Ь���4m=޵��b!38M��0]�������[���6���9����ED��3x&�o�4:�il3N(B@ȼ��ƇÎ�M�4$_Z(jɃǻ���4�̹}��Ú��cƳ9��Q�h���ǆ3?p=��2.o�}|�Cd9��go��t�즄ƛ� �g��P�m�E֛Kj�kЭ�����[��/GMu�d�z�6�3ۇsӴ�Az)!0�M�Si����s&a$%	8&���Y4(Q��P�(X��!!�2�Py�:��1n�M�
�� S>d�G;b!\vM	�p�V邩a�I�퇻+�	J�B4����>QY�2����x\������9�DF�f6��U�R�y�
əO�1C��D�'/C�����ʤ)ڈ�z;	f$���R��c���g���6���(4���߯{"9��l�y�n=�~Аc`�`�G���L	Fɱw�ނ7�IB�5�^*�Ē���#���L� X��_4Z0�0a����ϕh9�ЌP4g�MʶJ��M���1���Lm�5|ʎ�;Xq��tzA��~���O�C�$I�#��\�����=��j��΄qi�]�p��:E�$�q��fh��#�R�F�qL?q�{�<&	�Å��� �c��r Ys�/to�wN����.�,���B�o�7���!�E�{쒬@��%}������G�~��!j��P��~�cm�\�Y�e�0��ŧmc4���p߽c��ں;\w"�f�6eś��t�Xv%C�{�G=7�*9�rR���-AQV�GR�^FK�)Ƽ���V��`=`�	�7p�c_��Ϝ(#&&#@�_�y?m�p�F��{�� ��00��9g��D(�7���NV�F�i��20���4�d�2���pm�����ֱA�<�X�Va�n���]��/Zr�ÿ=m�_��_�N�D����14okI5�(�z[/��ۇ��oj�t��Ӈ�8�i8��C*+�05J��[$�EB-��C�t�,/�p��jxO}�>W��6�vP�cD�8;��lo�	��-�n%ĭV3N����ݿp�$a1j; ��
���',��wpt^��TN|�����oĝ�������!jl�s����AfeH�A�<tرEh��P!�f��)2�D/��pV��g�x�s�%
��cD�	bͼ�n���|��JǕG䆶�����?��FO�<o�K���R�����K�<2���M�΃$��6)S$��}P���D��WU��Lh�m�{��[�kGl����g:������T=�	��`6$�5�R3��M&�����)��C�>�U9�ǎP�oF�*4Ttn���cj(J+�6RO��ݗҹ��w�И�j\\,�]"�]�ݔ�I�����d���Ȣ1
r$�L!�@�i,E��А���QAD�#5�ɞbs~Lm���2���QHl�L6��:ӑ�Ǝ�2L�(sa<ņq��!h��V&;�𤶊;������N��V�l¤��R*Xo;��tÚ᭮���^52ɔ�䄅�ԫ�$$6`;���D2�	5"a��Ic��:@�Gw�x{���r����CC��0�,3�V�6�0]{�K�M�D80Ll�d��6�l~{޹z^{�4�[V@:�����W=���:{�d��g�7����QU�ù�'k��3p_]\�\�t��;��b�(b�q	F2n��35��g=���Ї�Y؆�%���i�#tt�+Y��t�݁�&���}�s��n�k�ק�����;U�$�bKqٻD���8���u�(���6���]�q<�s՛���͹xMs!���T{;�8��(��7��:�N�x�r�{����]�x�1]s[�+�TSȩ�����֑��BM*Z��n^5��v�]1��PE��9�� ��l�`3�ا}G�Q	�0j~����1f�DI�>$�:���k���VB2�B�it����O�Qa{j��/i��p�)&���vj'�1��^�Ա�W7^�/���6x���i�chH����3�CnN!�2e!��g��h[��k�o\�֗�qgO��8�
�y�C�/vD�1��V�w���;n3�N	e��P7xp?�p�E�[z�rΞO�.tal�}�
�:tS�M�l��,�,K`�9�=��?�h��ս��^:���i�=앙��W��q�Y��ۉ4��ϐ��N<�	�9G�A�:t�I��#
���^���4f����ė�3�]�;���X��E��:����Ė^m��C1�����9�q(�d��w�����զ�07q�C�ҫǏ�h���`��>X�*�oБ6K`�DU�gD��ɸ0���]\H�!=�B��3q��gfi�O����B�	���*��w+6�e��E�1ҭ��ZR�5]t��TG.$�d_uU��D��~���9J2"#f��UQ�R��1�F,��C�o�Ė:�f^�>qb�'���w���<��b�&��*������5@���,����8tftg{��>��l���az� ]�onZ%�@��h���\@��&�8�����!�N�5�{�%�2��6�&�3(D!��mϾۯz���		B�4�L��d4bQ����k�۔c{潧�������~J�*��������Y'�a}j��ς�8wo\S�U�J5�li�/[!��c~��_�(�ReO���}�°O~>��0�χ�`yq��/�/wb�G�w�7���8{��"PEH�`�\x|�}��g�9<j��7��x�(�W� �4x��������q䍡��鮎�8E�C �O�| ��Y�J���[�_sֻR�t661�Ȩ�+[��w#j�����6^%ӎފ�����n~>���]�b������VT$�������� �	:Vg�s�frV��;h�Up�퓰�x��x�&�S٧BT$7
����d�K�U[���������f/F��U0�"���ΘA�|7�bcm��m)ɻ�����`��.��-��>J%�V]���Pj��:'/H��CDݓ;}�V������H^$��A�n���b�!

I�$h� ����I�ܱ��6lݦK͢�r=`ƫS��d�v���:�xZa�@�a�A��ߤ����3�r��2��q����"�����Kp�� �h|��P[̜�hc�T+���5�;��+I"�E�ռV�svHf�w9�B�`腪�6Bi���P�A���v�DD����&܍����p!D���U�E��@�F⛎��X��a� p�'p9�Ojp,�p�Ae�	 p�-T��0��dI��"m;9�N���j���3Ib�iҎ1��z]!��#9!�K�|*Pر�b�7��������Kį�
/HH��p���=o���]m%��ɩ~���<�'�]�x�G3�Xr;<gJ�MWu;���*,��1{�����l�E5�f�i:��l��+HQ�%�bcY"ۦ�=��U�`�Y|����~~��\fb�T�C0��6]Ff�èmر�aVL؊џ 7	�+�!���$��)�-��M,]�<c�$��׺g:���"��o��QAv�a���K3�Y���"�ǐ�m�-���p\��2;G
F����7�ǆ�˦g�^Is�(Բo�s�}�/�H��F&P/4e�\�Wx܄�$���H���*����`tm���S�a��yq�˄ˇMa��1��Ѝ�:UN�Wu*��U,�8;���L,��v��Z�{n�u%��U��Lּ2o�.N�2t�E4�yn+O�&���4�'_*_H�ʽ��GM�Թ7�)��8��ꏍ����B��EX!"Q��l��)Z�&7ݿ���lv�����R��烯`�Iȶ�h�:7kPh�&��L-��M�\i�R潍�)�#�`uK�Y���4��hň�ƍM����K��d�.�������}�l����.v�z��
�����z��yC�]A���mI)�J�踤�6�)qG��L�c��w;imI�¥j*:�X,<�=��d���=V�|5������$�a� AEӽ?�~�^�6YOݘ��<��R���c�XhAUl�E8�9���5�UN(#j$P��8+��������]�nUېuM�g�8-6Л��:+Ġ��ׁ!o��m+]9Z�`���9�=�#����jA$��[&��˄��`܄oU7WC���M�c�(GI�	�6s�x�f������w�a�٥��@�~�`�<35�����p��ѡ��ۀ�m��Ruɣ�${I��1T�)������T,�әI'/o�����岧6�p����-��\8%%(���m0p����p�,v��pQh��$�I��Xʘ��C�b�뭧�/�����_��$3�=쐆��7Ѿq��y�npJ����3�5��x��٤�A�&8*ܽ��J3/8�� M'�Nu���ӥl�V�xi)p�-� Z1�'�ώ�a�,!�2����b r��uwYж��GR[:�i�84�p��;���6oTP��@�2�ι���q)���!-ȉ��j�^lG��E��I��hx����0��"�0��Gh�˼���px' �T%:�%	�|�v�(e�Ƿ/�%t]�U�2���R�@���H"�bBj�n
b�p0`-���p��č��=�� !3B���ϔ}�
!�N	�#���`��V0B'�t�b+ʬ�=�Y���H<�l7cbm���N�5��!\��O��DC��I���r3�;I[��ԽM�t�������Vy^��C�X ��l��r<�:�nh��Z��拜��zǰ6��n�M�Wdg�LX�Z�=\��x*�4Ѷ�S�e�-���>��Q��^�<1��/�v����S���é(�F*8u�_W�GR���
��l�m����v'*x$8���J)9�6{[�-�釐�a7tߌ��}%�eZk���&�H�0��$i���RK^98t�s�0]���w��|4q�4}�Sd˪�!�ժsB��J��28�U����O4n�&c�r�u԰Ӓl��1fǮ�Mq���f�X�t"��,Se�-���N��c�'�Z̭�>_j@�[����aXg�~�������`�29궓�����m�(m}x����s������r�I��9���A#L���Có�`�����jy�m�
�EӢ�w��*I%����=��E�9��꺦���U�)BA���.J��4�=�a-ǩ�>��e7��	X�a��\���oϯ8�B�+����l���b�G�����ŷ����������=T�$#�s�F68���GQ�T�<���XZ��"��k0cC3j#n*���oOD
�gvʊɰ��^�i�@��)<̗�$.���mU��@C��a�V_!�+��2-�i�RA!�1A}�R����On�����F�?n!x���O�M�� j��P�,u�|h����	/�h���֐҃<�e`�Y靁4��0�"x�F�c6��E�õlT��noc�VeN���;U�-���B�U����@��I��e�Ub��C>#٪��v7j2>��Y�sZ;���a^:h79[dl8��r,�\nA�D�8������-3D��uV�T)����B�b���r�I0z��]�Yӟa+	.W���^�뛺-m���s����7��?Q����REyDܯ&,�$�x�r[������{'M�b^7�Xj�l�Q��Vҽ3a��(w֐���cf�L�	 w��`.r!)ʠh��r�@w%]�B��n��$�H\�B���pH^i	o�@%�9B ���lHZٜ8f��jު����|�+�	u��q$i!s�$*$�ą=�Z@b�î�ѭ��̒�����{����y���k�S�^HK�_m �֘�hI-0I[I)����~��o�̮�9)�S+&�=��M$����F�X0Im��{@���t�.r$����;�:�/ Z� '9)#BG�B]<�x$i { %�%�,`(ė��X=,�����Id�*i"�{Y[�5w�n���g4�΀re^`%����������,|?���f�z\ɟK@�����]�Fv޾JǶ8JLRD���5�$U��4����!p�T���q�����5��c{���%����Xlj$YGKcbC�`�����Z�6�M����>�6���w���͑y�����Z=���L�(��ۺ���Y�L�a�{�!�G2��+��v�[9��Pls��4{�}�6�'Ci1�?����pnE�9�����;��\ҎD���P�P�p��;s0�h֜��:���[0Zn���d�,���]�r�#�����������|HR��f���GTj	����8RϷ�����zg��p>�)�+���R��qA��{�'���~غ�˳1u|tY�ᑇ�C�6B��h�;�i�:���=���$ѧ8�Pm��|2|y:^O���o3OZ�����{�N]���r��B�!����@M���"E3Q�C��(���0g�ߤ�ն����*�C
�bN�7���I�D�y7�~?LIdi6T��-��<WY�k�3y�m�Q60�l\��c��@� P��!��|�ce��͐��A�1��\>:E`x|f��ߙ_ECi���$z�$�钺�7���b:�^��u�QK�[q�W!j����b[ȿ��壿s����Yے��\vgc~3�u���z��o���0���(�{a�@��{�n]BJ���l�n�YQg|9ѥY:>Ы1{������40)��8Q�(�З+���?Z��X�f���׍!�B�$Ȝ���JF�0��.m�N2c�e��]��NJ���Ϳ^�����L6�b�����G���~+�#G�߹Cecq���Q�ֽ��D/s���m|61ͰM2��� �<h�o�Dz�F���.�*;,�(�
4v��kϝZ=z����͜k+e%X�R(��X�4o�u�q��b���3H����+�Qv���)qxD:у�(���ab��e��h/�C֎�n<�}��n�LW�G��D_}��p�a?��N����]���C��0�f"*���/�z��oT������ x��Vi�4F�[�s�k�"�1�YUіͽ�"�N��|L���Ѭ6ޡ!\$5�s���)�M��(�HƤ=��[�Y̬�+׹R�s���Y�X�64�<
�Cኟ5c�Ɇ'X>Y6�r%��x)xm?3�z�� �� M��b
����aTc�I$?T�2I#u�P�CHE�Y��T��	{K����I�u�B?ݗ���b+n8�k�#ƞ-�v��c*�7��e,�f�lvצMж��b�f��1�[h�i
@pݼ� ����6}s5�=�g!�#���q�8�'o䌏ɺ��"^�m<9�k�gf�<��$��yznM�@�qq�v���0X��kn5O���p�u�3���/��d{ m5Z���T��б��[�\>��N�ͩ�=`
xy�Qr�Ew9�`���ro�wC��OW��+���~u���p�$	C3%��I�W�v3��c�s]\�Þz7���~�,w��M�'��Fۈ�]&'�?��C����8<�?
�c�w	28Kg�b����7=�h�x�Ö�Kj����������K��+�/3��
���ݎ�ܲ�;�D4�n.w��?{��������l;��}8]��:�h�N_å��c4����p4�j�4z��ǟQ^Q��V���<����i���!f��.j�MݝK�y�fϢgTK�ٞ�m��[�����:6<h���G^Ƽ:7z=}����7�a]�!�=����g"���?4��Pβ�i�z�����|v�8Z��ǫ�>�+]<P[
XX��gŞ2p
Y��{3��>������3C���}���]%��a�Ʊ�a���;������3u8@Qz���jc�����Kư�'���C�/�p��ճ�+iC�3�k5\��T?��Vl���e�A�6��>��ܓ���u�oF7^ګ\*-�?P~�������i�Q"]kơL����2Ɩ��G
1�1Y_q_DD�ci�ހv��W��>G���A�����R�w2���*�����?�A�4M Y�"�'�#zP�˪�i�T��j+H���r��mC�}�������]�g�q5u;����o�U"���U�5]q���9��-u��O�.>����B�2�(Q��X|@��7�W�o��a��ND$&�P�A�Mm��ٚ�n���v8h7�a��ʺ����#�x?�6|���=�Ŧc0e�i����r6�����l���1Z><�z;��'���op;��y����5Ƕ{c�oz���������c~�|2��O�}���W��6ocsM%�����g݅��v��K`�����9�Ϙрt�/i��ϫ������Uu�i|u}�cT=0����H�0�������{ﵬ�%3RUڐc5]�wZΞ3�wN��Q؞e$k�L��n�=;����(�9B�&�ɖKl�7����gŝl���t��پE��Dmx{g7�xB����zD.!���o~O���w��~��,�f6c�].�� SZt�.z�3�e�A���H*�M�k�L��B�5�Z>�����nm��[dW��~��X"
�E�۫�ޒ=D#��JW�DᱣyM�zϋGk˝�&1��o�ꍶ��F����^j�ի#�y�0��5�����Pnv{�P���J(����3i���&���ʳJ��	�<m�!a֗2�ԞX�lll ��p�?`0�7�y�pS�	����X3�ln��ӻ�;y[e46�1��EDؗ0d�����6=���p�f�pg6y������xB�T���{�����B�6ݝIZS�����<Q�-�����x�MuF����ӑ�̞�Y���J,}��(� �tdG8t��tf�i�_�9�y|�i����u8������=	ˎ�ڹ��IL�B8�2�����m~��/�篟>Mcnl�b����у\���`������^��A
�4@ ��(^���l�Cmk|$+��{���]5*��
���>2ƻ��B/^���H�ʼ�O�������w��\P !����&G�^��7@�i��Ӈ�S&H�l�Ɂ�o��|���E��|5��8DQ�>A�4�^h�T����Y�o�š���dQ{��?v�������
@�Erg�y�6,�p0�		�����N=x�q.�X�iX�w�����B�c#5����f�{��MmR����i.�������-Mܣ�*�ʩq�+fq*��3�6�®�<�VC7���o7�{����k���xx񣣦�"w溜*U���WmA�tCK�G3����3B�#43|��ܘxغ�CYض8��|< X�}��[nW�L���%���AKh�0a�H��0��w$����L���6+WB�ܶ�g����c���}rk�7Q�5X}�J�"�_�2�ll`�6�E�}����Ɗ1���5gt�Z���՟X!�pe3Mb�w%\�*��Q%� m�B?��/�|h�a��׎9'����l���b^ lg�5�7�`����Т	���^�l��h�����٦">l��ců�E������ą^pʂ���0����i��Q�]��b�7�����/(�St�[I�<�qh}��M��~<V>���^{�n��)�v9z�Q^�؉�^�m���b+Ͻsc�%�4Fpa~��b<�9���x��xAW}��jSg�ay[t��φw�Nnʒ�*�q�wd0�H��#�Q�\��� ��Q�~��g��w�qEe(��DhɲB��i�R�F�����8�Q�*N�64����u��ijtU^yU=�����ﾧ��}\�bH�J{r⬌+���i]]S�g������ދ�0�=a�9MZ�
���#M�8Xs��$�ĭ��!�e��3<r�ɞ)�y�\c��޷-�ԛڈٶu��p��%��F׮[�sI��E��.�ǉ���w�G&�^�A�Q���)a��:�c���!�c؞4�g�>���̚9�v�d��W�s�֌V�b�Zü;�:1Σ\�p��Wi�/Cρ��؎s�A�l�����k���C�_�<�h�v,uT;��ݻ���-WwЃ����(�a ��f�w&Wg�O����~9�'���<�ci�}�v����5����-<7�����v�XxU����������� :�g���^�~�MG|���c7"Q���.�o��}��Ƹ���F2�YA�al�w]�߼��]�cnŒ%<�|�����7�tj�z������n#��e�!�����s��c5��?��`C�c�K�0���5�7W�}�G�у�����Q�!,�rU���;4u������i�����M[!z�� �m2���Tѷ[�,�����}�k�X42��8l���gGѤ]��9`c>F��{��:��T��7�7}�V�}�5u���G~n�)���kv8�'غ03�>�!Iu��_j��sL�_hج��O���^�&>�^�x����s�����u\u����T24�s��.�д�\�k_v����<��0h�KC�u���Z��:Y܈:�0�:�EV!��JA������}���Oelo�M�m�+��ҳ�!W�W#ؓv��fi��]v�r����w��[�+85�J,�:�m0�h�[���m��0�}#_{���݌��G�4S[n��1�ȗq�������u��u'�<N��}��|@lS�����M����)H�K"Q'�]-���D�b�q���.x2�a�į{�=���u��9�paӌ��06��ƬKc"�p�/���o2wf��?�^�=�
K�``�l�u�����ã�<�;�F�(҃a�.gzHNw3���5�9+F�m��R�:����޷�ǝ>(-�4piq��`VZcRF������{)�F��X�kГ]Qk�s��9^��ď�8�vۅ6���iovﾪ%�S*:��zv�/�kP,h浾�<x���|��_>��^eL7pT��åy��k�a���t�3c٨�ч��[�ulf�p�=Z��6,��o�%�SB]�2z��Ƣ|CМ/��P}�3ᤶ2��7�u�ͭA��#恌^�q9�&4M���n��:�H�I����%�з엷~{z=��c'�9����rQN�9-��y]���ڮ���7QV�Qi��ۉ�:��uJ$:/3�-�M%��It0���n�i�(��o��5�e���ޢr��,iw����6Pc,z'�~�hC����m�]v��C8��a�&��D�0>x����og^}������\4Di�<4}�[G2���"V1i1���,��Z^�c�V�хzy��oí����R����G #��C���)h�L=;��R�yguA��&(���*≂Q!%E.<�P����~9�@a�{SZ�����i�۞�%�d��%xl4.��ө�w"\��r+2F������Ԯ�D��=���S�ly���F���1�����lE�K�V�}�e�Q%;
+S0t�C6ΰ#>��ڞ,��٦ �+��P�X�߆���M���xZ����ma�R@����`�u��^��=��~���gR2�D�J����ґ�DPҶ#����w���G�ִ�X�봺���z�7J\D`Rt���
�4v�u��KJ�@�g;̕���I�$����E�wDڬ�N�h�9�1x� c��c::ɑ��M>y��͆���e!O�~�lM���n��C�[J�}��V�P�D���|h��:Ã�h/��(ϵ��oiG����y Ƹ�B�ȆD��r{�!T]\��i�����ձt�"ػ���dd�����Df��*����/�+ĺmF��c<5å���ǽ��\�K�F��Wj[��U�W�)ph�����9�BI$YǤ:�S���Rq��<C��EN7���/�k��ϵݚF����CK��0�c�u��c��/�/����yӹE�Ԓ4aI��^�ک�����܊�Fu��p)���c#�_L���Y� ����DW��}F8⡧G�P�{jzb<�+u������>ȝR��7��I=Փ2�ƺ/Lɬ�h�qЮu�Z{�.�:~_ ������`���͝��֥v�e3���Ą��ª��P!���2ڄ�N����C��6�d3��;gz����7ν{G
5&ƻdZ{�Y���9A�-�EQ�q����7��-[F�¡��۝%�k�xTm�#�٭�*�7br3;e�6݊^�f�En%��)
qS�%��f�3k�8��hu�.�&�B؍��͏[�YϏ��ǵ��JsK�lq�3�Bգ}����~���ͤ�H�󧈅�(�o���x~�[��0�8���Qz'���3D|��'_���r�`��x�����8��9/Z��uV�e˧VP��u-����H5f�5!ќ���e����.�\.[�w\��U��=3C������/���$������0�6�0T6��"�M�j���ɬ��kCl�#�Fn��w�7Z7n�)����>*���iJ�)�I��;`�;H@�ӣ�|
LAn!�-�C&��d��4����!~@��<�^��_sA0���c�&|?��Q���c�xJ0�}��w{��t���;���J�y�`\�^����g���OL�w�'o;nd���h�,~'�y��W��S�kB\�x�[�c�՛�s���C�.��h�^kp��K�]٬dn�h)����E�������>���n]�8�^+]���9��c�`�{,�U'�!A�rd�Ţ:�r�g��w`�^���Db�pg���j�6�('z��P��W��q.'��۵���ڴt`fί=L��,�Ul{���e�̖j1�I��ɘ��l\(��9�PWCɠT���g��s���?�/{�a�O����7�ft�㎫�|�f�v��yܷ&�:d���n�g%��&H�o&���7�*bT;�1ҫU|�b9ӳ��aY^�!�L�YͰU��;�z�5��Y��r��#�y>Xt.�����k�~��.��m�VA��+�����Q�[sVtD�(�d��]3��S�x����w1}�D�]'�y�,�vqt�����+�@�<�h�7,K��}�w�I�6o9�rJ�����bW��YY�Mb��=�t�ä���;uK�F�9UW�O8UmEL����y��fcH�4��}t���,��M=�&jX�ۖ��C��kވ�Sbѹ���V�b���)ɇ}�t	�;�ѷ��*|� ��[�����wv��i��'>�r7�@�!]��G�����^-�4?���]Ξ�[Y�ثf��Lv�)���Z�k�'���R}�;�۷	���QG��x�C�����U��D!�f5UfRkN�2~ݚſV�剝��Zq͓w;�q�����7��Ol�l<S���n+IH��Kvʅ�v.7�=Nmk6�-�&Nf�-΁�x���:s�vɉ�\9��G#E�����DI.a.�tt�T٢8&#��#+��j�5���tW&�^n���;��X[�\�3�tjChW���Xk���\�=`=e2	�&g�v\�.��
����HĳC%5���KuŮ�!�X���t����&�<��\v�ۯo$RH���	j���LrvM�z:㘝kC��L��Ӽ�]ѽZ��5qS���v	E��}>n�xħ3���{7
pB���8�v��T�N��!��0�;��ہ[�J��x�*�v��Sh�h0�"�c���� ��.7�u�*�Kq)iz�q]c��3q�c�n6uӷ*ج��!�L�&�ݘ�ԣSI�TtClv��r�h����8��ѹ�Z��@����]q�{Oe��6�e�P\zH>y�|�-_%jbY|�o"V�0�ugQ����iّ�r��ܦw[˝�Y�����{;��AΛ��6�N�ʴ��z9H]�]
,��Z۶�svE�۞�m���g<�&�>��,����y�	'<r�܋m�d!�9��u�5�p�z�<`+۞gځ��+"�FBU�ap�к�|j�9�*C7P���u��SG[2�X4&��2&Q5����Z�'=7#��6�*�ɵ�5�+��2�'P�)703�l�VÍ3���3�bY�q6�i�9o\�z\Se�v�Wg<�|�ۋvn[�w[��iVֻc�ۧf���W��C��<�ɒݔ�����;�Q��3�Pm�b��Q�&�N1^$y�d��.�ݡ73uĴ��]��\��g�ឝ��s+��^�7ۘY)�����X�kpT�KE���:��[��4D�[i�ZRԒ3�865�&�$Џ#�2�-�W=)r�K�\Vw��I;]�k�Y�^�S]J7�^�n�g;����9�^�ؗ�:{;��5��G7�c3��n�E̢�$iR�E�c��	a�nY����N�6�Y]�/����p�P/� E� +�$c[ m ��������]_!���\&R1�b
�i��YHu�!-pڤ���u��+�����/�؅LB�9IքM�*1Ԏ�2��@�q��!j�B4���u���U��̾�����`�i�E�"d@6�d������5��mFm����+�EU(S9��BI��r�����*�ci���lB`}D�vG��7�����̘!%�x*�R
i��D뀊�Ir8
����v�|�$y�kQ$�]��-j$�UW�� �Arv�q�28�WT ���q�;�%�%5�ZB޼��ʬ�;x�p{�'"8ėZK{� �%�{D�W�G7�e�e��R��̬��б���㘰�B��:}f��	�v��\���	T���]X�Cg����mƹև����Wv�Nr]=D����b�����v��x���Ұ\Q��*=�,&��W�3�r���5�2],rW�$y��;��r���jٸz�X2
=vp::�cN�m���vnK��Vl+-t�LZKR���y�lny}m��8�q�>�J�-�n]�?<����^�{��g 7G!)�����7Ʋ-�_]Z�ɝ���\l[gN��;/3{]���8F8}�󅐀���Ϩ��CZ��։�����v�j�M���/�k�v~�'x|��M2���x����+�p��Ǝn����v�f�ip�]��{<,y�>�z��@�8<j�!����CA+�;q׾�����Byk�I�l�Q���M�a�Jb8n����Һ]Ό�6�t�A��ǯ�ۿ�$(Q>�G��(�F3��ͻų���ƌÃ5�a\��85o�{�;��^J���F7��4��v{����ÉC�����Z�]�� �֎E�3�rf $	�7�Z�%�����������I_A"14�b0KD��	�|{�[[a�[6;)�.�w��1u+�Ć��2�q��Ye&�	Q���H��FQ_IB��X�!����I�m��LM.�v���2���I{8�V�3�bsp�E��!��O��0},̂(�)�d�(�5Ҝ�/�znaѮw��}�p!Z��xU}c(����e	����S��
���5ߦ�q�r���(�dp:~ ���C�(	4�|x.3���Zީ�)�K>�Z��nj�xY�ٗ�J�}%�]3����=��bI��3yK�����D{QA�) I=|$-DCb�����xS�3�KĈ(�����R��!�{[}������B�_��_rۢ�U.�9�n�Y�DG=q�s}�O��i�f�Yc_�/D��
�����'�>�Y���C�0�(��la�@���*��6(C���@��"0��}؊־�!r��r鸘�v�mZ�{p�퇾�7�q�t]���ፏ���D��>��j�p�#h��N��{�]{^�0��N5xB�g��vC37��צ<��l�I�e@�(���<Qpy@a� �6�L0�Yt�b6�ScI�b��nۣ��O���'��}~�f�ܺ�*�Zv��6�n8B���36Do���t):X[�>$(�\���F���YQ�=��Vdk\)�S�2B�_?���3s>�f6v��W ��c��8F$n��qZ.C��cc8T>�C�Z0J6�hol4󝯍�b�6^������T5_CC�Ǖt��6~&ΐ�|�q)^���Ȫ"5^���)�9��B<���특����70�Z�fN�� !zÎ���<���6��/��זf5>�7j� �،���!( q"R7=�n��lw��u�)��4�r�P~�(��?lZ(<O�z����^������uٖ�q)Fb��2랭]w�+�gH�ֈ�3��s�_��'Cae��J�I=�m�7s1G����"�i��)��p��T�z=�>���F�`��$p4Aத���d�d|�@�;��Y6Q�|H^��7�̄����\;����<]�����n�I�-��֔3��3ƍ��dwd��}�y�ǋ�y�jE	�7 ��I!��_�Ol�n�����>�����t{�޼O��ᝎ}��5nt��>�ݩj�!mĠ���EЀ�����ZE�z�,�r41�
�Hc�p��!��=��o�TW������	��]�^���m6�i����zN������ت~BA
� ��� t��B�H����7��,�[�+�6;e}�u���-2���}�;���1�zM&�}�i,[��Ī0)��]�l���3���B����#]>*Ǳ�����)�$M��.=|��=�E)I?m�t�
ApMd��_o��+P�+k�Αb��S3�b�U ��ǝ�PJ�VOZyF:����)�*�>6���ģR�wMV���ϢO��%�6z_=�<AB(�쏹Vw�f��U{��}*|j��n��s[�ϓXs�HR��d5�w��1�8o��|�|^��]�����y��%��ٴ��5\mZ�]ыn�u���Eg9���&����d�Ϸ۴��Mu79C������ˣ��{M�3��,-�[*jمUi�O����}��r�קz�S�V���^,���N`��M�
�����:,S�0�#�࡬^�M��D4��l\��.Q9W�h��S�yβ���w��Xw��5��h�CiLa�>(�!+�!},������K�{�=�b���� Q�����c�A/�����8�t���of�o�ֹ�z�~�F��.��O�{�m��B
��k��l"�0�(�`��0tI�e��;�Ǡ�ŎCʧ�$��9�R�C�����fC٩�⥜�oj��D�#��1�&�m���;/*i�Z-@@��'�X�H���~1鯸����j4Cy
=C�<���9���h����$6;��]17D�qD"��Ip�!�A��n��i������n�[��k���O������wJ�D�[v�����v�ۚ�(���Ln�|p$���m���>>��[Z�f.��Ch���a�+�\�ٻ�rڧ��rO��/EGqtrs�էO�vy����p;&�-���;L��ǀl��n1�Z��9�q:�[a���p��^���מz�Tm0�9�G���<��5�+�+�8�x�.��BڈW6Y�HVțc;FR�3\���鴉�o����'��_}I��JIs%ښ�d�G�Dmֈ���p��l�bD��M*AN��g�ɛ�7*]7.�A�k��=J����xp��d��Pq�@�n��*�ѡ����a��	
�"I(Փb��g��q,)�����z����{�����U��|u������6�4���zx�5	¨�B��f�Y������}a^"�W
�*�3��:�n۪j���z��ä:Q���e���{K=�l?pas�/�%�W�"�-"�U��}e�6X)�	��EPf�{�f�l���7�E�t�������xC9
���S���wi�ٲ�I����Z5���6�^��T��7lIs �!���Xw�{���G�wtŃ�4 ����	C�!�����HG���x&�%
E�|[�\�v{f�l�\ �e�V��.X�nR�ve��ՙbЈ�
�$8x!E�`C>��K$(d���|0���3�����Ї�v�x�D-i�K�q����r�6\C�������Gߧ�99<Ҩ�ȼ�6T�#��+����q}YAO�v@x���TF�l02P��z5�D��wJ�O��Dm��+&n��CoP+�[��v����kN1��y�{��M>7.4�W(Fոf���3.�3��>VW���hu�e���G��
�1�'�\,��Ak��e2b !�v$���$$0GeP�L1��M�j8 m1^�U�ر�׵���Cf�۝��T��X�
�nB2����\�=g4j>�	�fϰ����Tc�	�D�L3�ɤ���B0;������s��;�3M˶�Ӏ[��	l����A�����r+�XAY(ʶ{�<�����&�>��|�l�p����m���D?�A����
�Ĕ3�H���f��̫�']q�gZ�N`��t���?}�$82��0�S%�(�?�>�>�4!�����txe3t4hp�����[�h�Lf����R�wZS���WN������m�6�4������>�q�MG�!õu��,�mgY�7�B�a>�3F�{��^*$VC^:a��>�3������Ff��d�n ��(�]�惠��Pi_��Z�<GLm��Ξ4B��_7�"l:�{�([��x�d;(�)�Ą�vw]�{T��;ӵ��SuZ�wO&�\��^�M�ŹQ����J>��g�*<���⒪����)(M��@��x���x;�l^�޷*(s���>�ć������F|��넅�ᄆ�N-�,�|?�@g����{��)��dAPb��ã^=X:,���HjӚ���,���φY`Λ��B��b�x��܆�������>�䘌����ra$Tݬ3z;hѭ�:�:⧖�ϭ�����,�E��	�H@�
�#�N�4���U{"���}���C@�f���?ev���ސ�j�O,�%��C�o��~��_��Ɇ�i���<�~���Vt���4Q���i���ci�1�6���+`��pvC�CN�4��A�A�i�Pۡ��u��@#'����jR=���o�		8�p�
BM�0�(j���|ƊŠ��K��.�a��� Vu��.���	A		������l(� ,q ��!��,6:��FD�h��P�x� �D
�Q#h�ۅ�W"��x4�ۇq�˄;�RY ��~�5׺�	�����"���Б�wS�=��VF�ʈB�m�ק���]~d@�0����eZ�I�5O�#vle��^�S&B�<4 ��^�p��0T�&�#���`���]���jq���>�N���E��!Y�b�'r�u��:g���n��F3]�p����V��f�nղ���u��e�j�e.g�>����7��L$��U]>�	C��y�����L�t�c��몌�ɐ�?W�rl�5�n��O�U��{�m��S(D��~����Wv���[r�3�3�5�YF}�c1����5΋H�,n�é�0	�/1�NpH?�w>��I��Q�o4������Yh$4o�?SM1D�Z.;��t3ۺ0�;���������X�I�4J
�*��"�܅i�@�J���B�)�	2��m������9ٟ_�8@�x5lil�+�dFd62�c��r���J��ϗ��@45�as!�[��JV�,a����h{{m�0���%n���^WY�Ee"���\�f�Ǻa��3���X��n2�d���x~B?_!D|c��PF�Ô���|�o�߯C��i�G۶S�':����2񃦸�l���Fޖ3w @�>q�g9a��	X�lik��3��=\�Nn��Vf+%����JXdƅ�k�s���O>H�SY6N�����ۥ�n.YG���3���m^��ـ�S���6�,�{�=��o'$63���9��)��w\��lۥ��,p�\I;�15�cf��d��I$��j����SZ�7+�}���;ڸǔչweĈhp����g8����'��ó��cHR_.�2F�bD�,d䶘�1��7Svy�9P�gv6-�/b\�Ѹ��m[��H0"��sF�P��r8��t8~#E����ƈa>!���|:<3�C�|uYgʠA��clk�O<dx�eW��.͠�,��7������"�ӡ{�	��0�4�(���!���{'V	��C�"��;�7�y�e���V���o�K7A)�@n�8j%$���o��=�z��A���p�_{�'W���b״�{�wg:d&�S]"�c �r�!�>�e����ڞ{�W�[c$(�͞c=����õ�}��B�<P���9L�ϭ�G,����x��
Q���
R�#�h�_ՠ�J�V�~)���P����:b�A����=z����q��w�ʉ� �e��id0d�.�3�!������?T���g�u�N@:�cq�tYn��eհuh���x���L�`T�|:|C볪��1�92�c�a���$����{
����y�oU�)��$\:Yl��0:��R$&a����	K�!"�QV��U�#o����r�̂u�ri�ZF��b�w��>����O��E#��}�߽�A��M{b�2%w��b��߲��ogOQ���������c�#�� hAq_X(z��M�� �3���i�h& ��yj.j��!f���M��뢗}�4lKW���Cl$&r����GN��� �$0�
��������`�1��&�}����4U����G�j�c�>�T��:�J��f�@�Dh�׺`��h�:dP�#���vX�9,wZd"�4s��2;F�aFҵ��v�����m�}p�d��HT HС�w�A�� �? 5���G��1����P[��t�ؗ�睊��e����U8yu�|������^Mŵ�!P���(�8a2{��=d�agO�
�M�fM��C`�ؘ�m1�Ɍ��H��;��5�޶�2� ~��8��ః�"�A������(��^/fC�v{c��������-A�������������=}9ag�B�C��8�7}8��Cj��uq�Vw�	��m�D��Q���UT)h;O�(�	2��|Y�uؼf̈́��Q1I��nk�fn-)���*�*o}��dY��W�k
f���R�M���O���T/�[�n���]L�IFo��-G���� U�R�{oQkO��q�N^qG�κ����/YZX�vόиO{f�Gj���Lˬ�n�b��"�`���vH�m�f�SS� aS�kk/�kj[��O�^I��Bu�d��&�v�3M��؉���͔w��3J��7y�7w�S����FLT��n�MUu�ݩU��,�Wf�QU}َ�\F���`�j�8%u���oN�kߍ�z��jBκ�5�1��ޙ���6�f�ˇ�����3p���l+N���5r�]*�u��fZ/L_NX;��]�wթQ�c�̉.P����5�о�)�ϣ�s��}��Խγ]�.����䥜9«���v�-��e�Fajm�d�&Q���Dtֻ�<�U'r��k\�Org��=�#]|wV���إ4����;��ɒN��ZM���gM8��"*���:f����K�{;�J���b��!�:Tg%�C)�w�=�L�ޚ�5Od��a�lm���̳?'�q�R�S�˛o���	fm���`5�P���V�X-B����,^���]��Cg5�e(=f@"��"_]�Sۃs1 �@����ڒ�B�i�Am�[�IA���~��p@kԅ�nRFw��W�r�F%;��D(h{]���槹��˚�F4�ްG4#5ܴ#��K 砯��]�3�堻�Y��7U|׶�.!U�����T��P�@޵�� =؃��Y\����|�5]�i��zS��8�l�<����
��ǭh�ѓ1�o=���b0�G�m���/w) ��@�T.0S�f�C�u�RQ.�a�eݏ����V�쀴ў��r�)ȉ fv�{7�z�7ݢ����A�e�'2���UY�a�1��ov���8�ve7�@K�wQ ��+FC\���w^��.��/x�ӷB(��\`��5Ȕ���9Sy�.�b�Y횻��C�}y|�؁�4BճC< �n4��U4j�Oն�@I2XCR[G;���)�4S|!�����|8��F�\,���`�1=sd^_�@0D���~W�5��r.1�UP��_b��WޢC�[kg|��p�ϵ���J���7������Ǌ<hz�cm]]��Ã_(����������X���Y,�X������]ԏf������\[�HͿm�����et�v\'م����0���Ō�|stoct�Z��:�4�ݳ�qWO�?O��(�	�]��""��%���	�;��x0H�6�ӞH�D�)�0�������"���+����'q��p�4�w��"�
$7��
C����̌c�a���AT�f�B+�J/�&�ra�8c����|����)�s��)g������{!Ë����
��K����N�4�gb2�z�{�#��\rIq�ء!�}OA��A��RGh��d�	+	���ڝ���<P��R����R=>�M�0_�eEGL���W�J��4A|��pw��]�OJ͎��̞ͱ4����os�׳ �]���}pCP���ԯ�Ow�y�/�i�l�hxv���:Ń��S �O�;�4�ne�K5���~��?��xCw��R�c��ݞ�t!�M�/�w�L_�)3d����f�x���i��6i?�ǿ�'/����$5��s�3��ÊQd�%�lF���(�J�.��T�JM���o=��ܒ��Hߏ���M�_�@���G�$yx��";A/~��#��#��!vl7�z�h�cD�~�}�H;����V�T�%���Q�ć���&;&�;Wo���sMr���p���Xhk�x�-�lj����JC0
#ݽ���S�m�To��� ��x�bB#�1��#�$=kF��?���a���
%�OX|�m�X������e��{�w�J���L�]_;�V����hB{��_���O�^���w�7�3���w���衔pg0��m6�.���e�wV��;UN�K�B��~��e���8��9׽���DQ{�f�ݡ��wą�H[�a3��q�J?RCL�p�'�� �
t%-�'+*�Em�uv.��l:��0.���T�	H�O��V:#��HCMK*�t6�o�� ���m���0�o=ڽ����a {�v�������۳۵qÌD�#����q�h�����2,e6��6�r��2c�qcǞ�n�+����O��N��Dl�<j���nz.)����vj��q9��x�O�ml�pC��r4��SIjjX�t��j�}պ\�Cz�Iu��~���Y�6�."G�uuуcG��Z�����.sc��rtT�P��	=p��f5�#5�K���֨��n���8�n�[��z����߹��M�,��~2�s����>9�Fn�a^�a����fowat��L��m�{h�ίY��/�+��!������\Q�t�%��<����G;d�z�8�"��a֘2��Q���|H��g�!'�F<��G�������8�n,��ؿ{�,C@��� 7^>(��9�WD����@��Ci���p]��,!��{p�)����Ԓ�33Eo|s|���y3���^%����j�P ME@��Վ�/_ӫ^�B���ϥ��=���Yl�R܎�����O|l�AC	��b��@��G�~T	Ν_��5�Nu�l�{���͡�r�ȏ~�Py��}�����H���y�.�f��]�u��:�����^zq��9r�I�F��"r�~ݙ�\�v���Y��O��/ �^��G�����:�4��W��ױ�o8!�C4�(X�dp �O(��P���N�a�8��z�>$(`?a�"�@��&����H5ե7޷P�+̬��~��0����!����A{0Q�����p����gn�����5z&$c��0oxh�!��&��_\��P�b� ǡ!!�/���x0f�_�W��`cnfDI���8�SE�BHG��+xxXB���T����/^�Ʀ�YL�U��t�2Z��g��e���Qf��~�zQA�p,�a 4j�!�p�|)�ض�Z����k����A�B���|�4=�u��F������p�̈́��l꿣��I�>*6N����~,�k�m�7w�G��ߋ���6H���̣��
:x�U�3��I*J"��i�7��$��(~���v��Nm���a�.e�$�bi%��b��ۓ����&n-�d�����%Ge�������p�o�$2�:B'�},�r��uȈ,��V{����悱�ý��BJ&���/l6��l�����=���#�}<�Ha ��E̊n$�^r�������G�}�h�������<���F��C\�s}&�@�B	���7۲S�n�.�
���j��.�= z������"�$1�����M���ԐnN�믏������U7vz�;�	��6�i.�uQ�*�Z�u���&8�re����cF�JRPP'�C��w\3�m
�f��h�]�]��=�=|2BR_���(����7�7EU8��䐤�p6�(#@��ni�	({�� �����C��e��!j��AxN�k6����@c�L`�u{
P�08��?@����H�{�7�
�尋�o8$y}�B=����Xn*2��
��2�\z0��¢�!��&Ͼ����Y�G�#k�8e2���d2���Wn��َ�-5�k��4��lY��	2�D�B�-۸��	�ßBT(�FS��g||a��8R�Mݝc$�tg��gawo��ز�~(e�k��-���]�J�r���j�"��_e�b���VQ�1����ZK �c��HQ�bf�����!vj�n��^a1���n��؂�@n˲�,t3��3�<h�F� [M�)#L4H�,�&|��\�Zs�zN���xD�(?)��:ވf ��
�{�}v;��%���)�E���+���=��5 y|�:!���Z(�,v���Ɵ�xu5P�c=�64��`���.��$pK��p��,�ݴ&3&x@X7�{-A������z��.n��Q��	��n�r�O������d�Zl���!��1���K��� C3[08Gf@��P�@X���]c���4@�4��Cm�m��gzkC�kgO�����<�/��I����I���b��i�b�\��[�%�m�/G<r [tV��o֘q	CXAd����Z �<0!��>�(B���/�U(��+ƊOM����9~7�*Q��v<3�x������2��K�!*��H`��$w~����8g���9�7�`62ȵ���^��K}Fz�A�-4+�9E8� ��2�!�$���Y���g�a����#z�L՜��r�<WŒ�2ІR2!Hш>��-���-���Hic����8���=7���aR 5Lk��u��A�=ߎ���n��������  @ΡZ�4d�a\Й�s�[A��ވV4ȥ�ͽ3lT��Ws��#8oYcU�!�)�tn�R�Lbl�)��Z��:=���MS9�A
(�!AI&�C�_c��fTK�q)�r�X���j�W��eP �\gT?��'���x�2��i��#'4�3��Xy�x7-uuvz��%��F�l�xM�������vJ�zw&�ɗ��磄��-9��<i�GT�����M��`�=��t�=�V�@�ەp䷣aK���B��=�c�uv5�r/�k��ۭ�A���@`	��8������y�z�<C���Xg�:�����<2�G`��m�U�[�u�g�UTm��'p!1x6\;����*k�!�\W!�����c��D3nlv���n�l�&s���a���s�nn�6��x�?(N�R��>�D��3t���V�$�5} ���c��A��~��z�Jd��|��~:Y��@l���_�[6clk�>������x:�=֮>�s����H�\)N@�|C�͎Z,��K��������ڇ���S����"�^�1:O�m�.G9<�4���Z!l��Hnk��{�ַ�ćŌ,�P"Bzg�a �D�Bo�����p&`1b�=���i����7:P�#Ζh��8����3#��A�晢w��l�8ZQh�>��O)r��]܉�,��հ�Ћ�
4��vm1�uCq����ǚ�����ף�ֆ�SI�6�I��,����?�U�3g�^�X��
���D������/fk��l��܇fl�Uў�����8�dl��l�r�"1��
xh ���#,r����U'�W�n��3��0gY��d z!��tg�7/�������?&-qO��~����tb�2����/��ț��U��,V.�[�h�zv<~�����A��LN}<��b抨7�Y�D������1F �Q%o9NrA��lTT�N.ٽP�� E�,P�%����B�}p5}��$4Zd��2r���
ʃl����#�U���]ʪ����TN�ݪ��у��Xt׌9�n���5��6>x��01����$!x!�,�	��p\B�aA�4�~b�iXϤR(�b�����Z�� ����^�͐�	f�80`�pH0�/��,\#�P�(wm:�Ha�sDvhd���j�x�\�
�𼧷��n���l����"ρ���N�y�2�o��T��1>�=�T;�Y��g�댯N��5^(p�Z�#ga�)I�E�X�;bm924!r7>l��Ǧ��gɰS*H�_��m�>ţd^٪��)S�E�7C:t����K��e7��r�����K�E��H���GFߠ�C�.>�b%Ą�&1̀���.�^�}k�wF�40�Q��Q�f������}��:cZ�x�5�m�c������������0�Z���0k����tj������ P<���m���/����H�U��lm�p��"�E�4�d#���$Y�`I|H�z���u�&�|%,#z2��� A$3�N�e���S�"��|�Nٰ�_l�.lp�x���o�������fzj����ԩN\�CZ��XK־���?��Et3�8Q���`��pv����F�[�ܑ`P��cc��]`�1�?�{��y
K��?]�a��d�&kH�z��t��7�i��M�ƛ�D�������'����?J|�)GI��u��'ǋ<�/V��+���@�&��˾y����8��8l2��]s���n�z�1�vK����M�X��ɘ賷jn"�y�k��؋)��Г������B{�+(al=��唬�;;G><5׽�"�YG������������zT���ԖI�������)w��@�Fl]?zD�����IOj$8V�Bٵ:Yj��
�{#m���T*!�������7r�rz1�=�s���e!r�Q�=����g}M�� �#�pBi������z,!}����|�~�ό�25�'|h�]��7P(o��	TD6���0��/C�]��dP�������QB4��g;᫳�\���ߙ\g!�M���-Y��/94�n"�yq N
�:�w� ����#}��&o��~�K�5TE��6�d�⑄�dR��o�N],ʄI�z�K$V�K&���0W�c���}�s�Bl&X9c�s��MtҖ���^n��])P�l<�m4��4���Km�7[��C�c��*�8Yl��h�OϽU�
�;�)=��0���	��AN�O]���Mr��6�t�:�O<p��)A�l�㒿j��jӀ4`2
�%0}�G]����J�ϊ�6Pa�Mhp�~ڦ���N�X��F�u�������P������keȓ�!�ݎ(�T��]|v2U��&}��иQ^�!n�4���8Ry�g��h��P=5��-4�N	$���A|Cg���i�/���BP��WoNp��a��r�Q��g�b���ͻ���׭�Yc�n�㭢Da�^��nٱ�tæY~Z�c*�8�����Ć�3�CRm��,���pi@T_���`r?3I�Q��l*P���ݔuYĊn��hf����|Y}.Ru���^��k�YGv8pfk�Y��{v�7���Cx���΁��������鎸��W>���L�y��{��$v�rMD�J�a��דbА!Y&*ǣԕ����g��EΣ��.���BD\�$�<t�4��`pq��~�h]��['`���LI��q�|�l8]ۧ�r���T��z�YT���hD:ީ}cI�g��uy���NCJ�e^5�P�u��&�Z�Լ��p")q�v�&i�r�O�-�Vf��wm���W��H����;t�����ۈ�w��l.{vf,EM k����eD�7�Ԋ���.q�xA��:����'\G_�S���]�b�#9��<^�l�ka0��]��g�t��{rjV�]��$�k^�G�[��Z���1|3�˗P����\��96:o6�H�1L�������'��r-�u�M��Ni������WՋ(VȬH�6(Őڨ�D�L��措n��qmKB�_2�F�0��ؒ<p��`�\N*R�]<�)�Q�e�v�ѫ�]�}v��6R�~L�ę�o���"�UR���7�)�8#����֐S�DcV~�D��/���K{ؤ�Q��r�,���j��}�qEM}�H7��][W�Χ��G*m����n�0FF1���6�4�?22c�U�Fr|�'	�F���dC��>��~l�8��z��'�n��jJd� t��g�HV/��oi;()R�Tuak�@0�]E����b�v��&�Eͭ�4Wp����1ěˎgp��"���i�ϸᴻ��f�Ĥ#�"E�g�/�w�1D2������J�?Kȳ�o���JV֖V2����֘C59�M��<;��iKY�A|�D%%Ժؖ��UC�4b�A�[�����v8K�{�ӝ1��F�xƞ8�ܹ;{<���e#�c8�J�!����+;2˪�M��p���
�<qq	��1����Q�D��Ƿ��C��.;2�)�!!TŴ����1�����.�SǴ�j랺�E�џ5�Z��Y�v��j�t�!����tkI�V]S���7gb��NK�La�NC���6�黬��yx����|�q�moG����c��CHs�x��r=�
�n+�c
�ݪ��9��*��e�Y���׏H
�f���8�� &�D�ٺ�����0n�h�}�iLf��v�!G;R�7�ٹ�K�x�'G/eJ5ӽ��vx���t��{���[�K�'�7��<v)�l�d��6ɉ��d0�TŶ�m��]c�n��G7%�p�gRKLk�d�׫:c��ɇ����n�3`����B덶�:u��L�ۊ�:q��8�G�m"�]Eg�i��A� {mn݊��nxn���k��ê�wQ��7]��C&�:���=B��ç>N�qv͉���r�Զ��.n��A�Qq�6P��m����vN��Z�c�zҏ���5�Jb��ۺ�8�K�����¤�]���@�rn�f�z ��N�ݍf��9����NG�z,�d��1L3��rFݑ���ڛ״��'A�`-k�ɽ�cص�ܓ�ޞ꺎Ď�BS�s���Ӹ��53�v��0�-v�+��ױ�1K�<�\�3��튴n��{`�.�joV�=z;n��9�[����e�|ʜn�6�0�v�6T:�@y�+�v+d�Tm�ގ!ݢw6[���G��ey4�p=����+�l�v�<b:Uv��zG2����6�6OC���c�8��Sg=Wlʜ���=�xG�Q��c۝�K�vnR�ฏtm��s<N,�N��jg��۫����3�����e{n�q==r˖�Y���u��ݯ4v�)�-kq���":\u�Yd{��kZ�]�h(h������y��5[�{5�e:�^u.�o�/c� �_4�'y�B�D���G�`��m���n��]TJ�1�Z��{P[�@��I�# ]��`dT�5D�_K�鋬W� �Dq��iF�\��j�n*��߮�$�&�~�w��i�����E���G���K7�Jk"ة�ح��ֵ�y�hɜ��kށ�7�
I��>վ��j�{��WǊ��Eպs];�o)�^�%�6��[=��݉�3%��9'�ty{��0��R�K.���b+�ez��vNTl�7zu)�%U�I9]���	D����Ȇ{e^�*��p�nln�6��3=pn/Y�:$1��%��H��s�LlB�EۯSp��5���O���r[��\m�u��ˍ��v�셂�x��*��Ɂ���n�ٜ[�K�(L���6�{'.F��ON���xR��ڮj�b4�$��Y7��8�n-Ovۃ(��6��.�p=O��C�G�-R��zf-Џ�;���!�m��ѻ=I��ܣ
�q��Q��7d��N{'V�c��[t9�,�!�Q�|�'a����(�>1@Ĵ��J�c��c� �/�v8!#c�7�K<9	O�{ȡ u�<����pˈ��)q �� Bo��}9��w����|(��L(���љ��`�_�,x\�"�)cpM�����z��z�:�C��\m3>DÁ�A׵��O��z">��]�R�9�-Md�I�*c��!�L���H}F>��{�O���p�(LHlw,�W����ʪ�+�cp�vR����(f��>,ћ��M41�+�8��"��s�;��gXz��FQ�i�#�j{/;s���s��bOs�ǿo�	�v���w��_s+�2��.�Bc�d��x�A�����H��#\��6�Ǧ��	b�c$�WM#�]�5�*)g!��Շ����=��u�>��j8�p���Z�^6��y��^$,�ڛً�=�f�Q����s�_o�`פ��{3,���t@�>�gt8R�1�$�,�����es���8��o��c|�ԋ��%SH�Y�|{
>��3���l�"��u�h�У�^���F�9��M�F��i�&8���K1S"�BZ|f��I�ڡ�ߋ�ɬ�^[�sZo}:}�Co��ؕ׈|�لDg�T
���1��^�`���SzppߗƩ�©�hB��e�/�Xz�H��?Oх<��Q��!BB>�U��|)lDV�!��p����,e����te�W�sq����$�>I�[+ln�� �Z���_W:��ηŦ��{�Ő����qx�۳H���g����`ת�æ��鲺�1�-��u�0�M��ۺ�N��og[����]ωpf�ӭ��GI�Z� w"����Q�:�s�Mk���1}�W����ߞ0딞Z�������6+��	��Զ:j��1E��y��}?G�v��#���gB�c�*=v�cѳ�G6A���FR ��=�b�0C3b��)St��Þ��M|R�(5����bp#r�g��^�_�P#(�-1w�c-J�^���u�2�$)4ovW��!aC9�G�Ö��~�Ah7x8�m��b-��bH���( 1�����yC �8�؈�(��b(ϙ���������Ļۓ���2���4�eE3=��̂n�w�����'N˚识��?]���J�������S�����l/}oD�9q���F}ݷ�>���ӑw�e�z*	��}�wur��U�E�,dDfĹ��7B[�M*�}�M%�|+�3�����Ć�`�ª�T���I���'G�.�Z�;�#x�ڀ��]A�@�6!sT7��	j۪��q��>YCUϾo���RO_w�/�4}$<��C�<C��[����"��b��j�fy��G�"���NN>������T�r$et���Yj����ҎcfHj4]1���Vh�D���d\w%]�H�8Y豚>/��-Dه�[������;�@����ah��� �.�A"B@Z@���G��1�rEI����uA>^@��
" k���忏���D^]Y������Ex\������ȰY�	2�_D��oD=����o�����}N���ˎN�����<5�4�׆��.>(�w�;�vꓶ;��1�{���2WmZ�/�[��ʸ�8,$*�0�����(�(���"Z�o�5��i@kh���HZ�Cň>	^$3qx�PG�I��`�rѤC�YbU������{9C��C��\/�w:��W�j�3����u5ϩ��t�9��F����� �&W�x/��?�|��$PH�*�I��`?F�GRU ���u�b���
��1��盿s�C�@ޛt�Ss�8j �}�&�L���,�� �ӈ=O\Lq�6�5Ψ�m�:â�cIj�b51���uN�u���<�A�� 
E�Ն�Ώ�C�-H=����o���>{Cvtfjá�����^޾���ZM.ؖ���7{V>T��y�!�~�}��]��v�5�����'��>�v�b)t`a�������ݐtr�ǣMt�D�F��$Wh���{�$1qaT<݋�x�Ֆ{���-�(�f�#c5��гcP����z��ꛅ����{i��{�fp�wW�o�,��V�l��8?�ةD�m�������*z�Ɣi}ʨ�M��G���5^�l��5^!V�Qq�rA��.>����ȡ_&ll."�YJ;�$:P����g�C�l�i���˦�RB��I�����}�|�!Y�?~�K��a���+�T%+�,���7�	x^-6���c��$�`+5Ĺ���v �B����W��J<2pϓ��s�IϮZz��i�Rnm�y(�m �$m]�z�^�#��]�Z��uҮ���C��%dZ�n7�٬sn�Kw6�=���:�r�Z����mV^����y��6f7M��+��f��.�U�1���#���{��ܼ�n�2!�t]pcm�R��;Aہ�W3���&:��=z^��q�2�8v�����{�.z��Mg�hm�\37BI���w����5R�8A�H��E�	e"K���a�w$o1M�2��i��;[1#n�ߕ�}�h�f��p�ߡ����7	�ga��Y�f�xc�����L��><�%!Ґr:(�c���ӻ��]�T,����z�Q��7�x�{^�^f���!j�������I
.B��k7��w����9ú���v�lۈ��A�|(XR�όۊ��~,�<�7�f������>��X}��vƎ�d���E{�~�喱��}C)���aG��#`���v��s_&N�uχ�ld3���^ET�~<6����>��O�l��,�f�霷f����	�{�}�ո���K������[�����5\�l��QF��d> F:�4��a��>����X�'�AQ�L��]�C��RQ�l&I,]���}*$q��Q�.N���kz\�i��Y�Q�g׽����B�۳-������|>� �C��%j�O��ӕ�'9�<|����&!�KV�HV<�A@��޾.
jN!7D,X�G�������oɌm�����T� ���x�B$,\�Y�6geޫ��	��^TU��fR�2���tE���p�79\��nZ����ʲL���9��E�Dt� ��h���~��r�#;�7�-t�����Qp<�����˱ʻ�VC�3{4���D���WP�!&��X|B�p��im�r�y�r����x�������|w��L�#%0mt$=��U5�VCwl����hh��/j����Da�P��<��&��Ho>�֊jx{��N�͗�6�8�60 ��xs�e8CI�PL(z�������~����vp�~4?��i�)z-у�`���}!���E`��`�N �D@�5�	��a0�|@�&e9����+�i"�����]�+����nɮ���|��{���K�K.Z�C�w�\�"�E��Å33
5ӆ�Z�VL������ɶ/���9qwU�׃t1��.<���{7�<�ߣ�..�9f��Q�rLeW��a������Æ(������.Kg	�!lC[챬8�Az�u�esl�v�Z�e�+�f��F����>��Y�h�"@ap'f�ɺ���mlW��9u�b�l�<rl!�XUɟJ?���3�{5�;M����D�=�C4h�PE?��̋c�. �7C����wfUܧSva$i�m�|U1��o��W��ѓ����og���^��wݍ��<�l���ZL~�.�V���������� {6{�Q�P�BU��t�K�]s�|Hh��	�5t���߉ן1��83��ŮwT<6�A�pv��B�f�z	\�8;U.{;F��]�z��E�X�ڸ����N�7(�j���>fsT5W^y��?���������ݐ���0~$�'�Jbwz���߫��x1QQ_&���g�q�jz��U\��d���A᫺��k��.��_w&>�g��$79���2��,��/�����u؜(X!}��=`�T��%QP񝔬��՝3�/�R�
���Jf�O�]�,�q)O4�g�A7��wd��)�����yF&�H����	n.ٰ��*>Piy����hM��ٺ�����{��(�=je�8l�YK�Y!e�<>m���m����g��$|H��ǵ�*/�!B��I��6n]�;�$��\7������J��۫B�`MFdMK���3�`L
�r�P�!*:�f����<��>�ϕ��3�f��K%ԷVQ.?�p���	R�'<��h���J�J����������<b����>���CA��l{3�8{b�������A�(8"J3���u<ix!zwa;<�hӯ�ޭ���;O�%��+�.{��UYM���Ȗ&s}nl���k�Ûhm&�eQ���"��$/{�¨�7�>��	\	��'�[e�ۀ�6c>�Ĉ} � �����($�|7���c�E�7�[p�m�M63kT8w�7�*���|}/�b$SvFT&��@��b���+ǋ0����ƶ};��ښ���z���X( sB$74H��li6]���=�t�neR�0�>�%={DDDE=�~Q���4���:��ú�l�ȵㅞ1��V:��0ÿv��^림$HBzp�9ƍY|CpSi�pvPփ�4Ɛ��M��8Z�v�~c���o�jnCz6,� �ч|��Y�aҔ3�k�r��6���O����	�-B)O�bm5���m..R�쿴�-�:�SU.�#\J|��xi"�we[W���?�a��z]��ͮ��X��y�kY)k�%�LK՘�1�!�n�#;�O;���n0&aq'Q���5Ě\E�%n]��ur�=�<�r������T�c����P�欮Xy㭮����.X�#��5�M��CB�6iG[�7la�㵳�edl$Օ�h͙h���7��Fފ�A�}[��'5�4u�X�Tީh��X�a��l���Ǳ���~+����s��^��OR�)wD�G�. �%�d�����wAK�+{QĘ"���a6��\Q�P{s2�C2ٮ%���B�ORq�����첈�&�i[(�D�/�<j����\,��G4s��ߏ�>,�o�,s�Ё��y���߸�ٗe��V���~�5��H��&1;�c��:���ӋA��F��Q��E{v��K}�](�0w��uo���Y(�LE'E��;�����"�˻ؗ�>$E;$��������W���:3[z�k�����؁��3��	G���4ޔM�L8*n���o~7�Ϭѡ����-|C�B��O�al��8C�D�ϙgxV�0,�0��'����;"�a�f'��������H�w(!¸|ku�.{z9��"��1�����XAW��9�½�������/�<��:5�ױ6':�ZmTnN8^[��ڼ��P[�� ��A�y���g�U/!������p�IvƆ8���6B͜���x<����G	����ߏZ�� Hq^��!�Roy����m��&pX��4��H?�h��Ey:��u����4q�xx�$y�UTn�KWH,��.<��{uz�S�d�y�{Cv���,y�0�������Ət��oڳmh�3}8j}���!��s�aH
q�e�@��e@~ps��=R�uZ$0Gp�����M��1����}Y�r|�3��#�67����6��sp��^����NPZ��1�.x.|�v����٭�o��\���e�1k�ޑ	hH {h��ۏxwD�/�MALR�y�o�=*ˢS�Վ�Y�Ҁ�h`�D��P�O=����"�P��p{�����������@xWvED��og�L��80���I1�t�bezݝ���j�=�q*Eñ֕�C�Yy������uc���H��Xʄv�k�g�����E�s���F��{��>�=x��i�:D���@5!�t�{�&�) Qa�ݡ�%s��Y��+���[�GԾ70�#�6(�#����CH�_}��03�ϴT�e�X���I1�~˒���캼,�-5eCE��=�ư�[�����h"F��;D����+2�q�I�>F�Wk_mR�(�ݫ���������C"
q���BDgh��5��ĳJ�^
����������s�w'><���:�oV��cq6��'"��,=�A�ɂn,ܺ�*��E�%T��ĚqO���]��������}�D�Fb��	B�Z���hO�$���t� ��D���EJk�g�,	r`'C ���bm(�[M͌����;r�O�"cng'X�D��Stu3�$��p�c[Q�$Lb-N�D�م��C�b7͎���HMl�	N*T��`�"v,�p����wRsr��V�Q)�=��h�QJ�s�ݸl�ϩ�&N�0���]����i�I�ԭQFx����̻�Y�|���I@n�T9ծ����ad��1��;LP���"���â���U8�� ��j,���s54-�p�l9;�ð��u�r�?(u���E����˴{b��"LW\}�,��>���pguFu�T,"�r��f�tlN<�/�0���k��3v���Զ�������F���Z��Y/�w@b�;<i�[��̆� 讁f�/�*sD(�^���_�R"�?�?l�ug����SQ7ȟ��"NcU��O�$��`GK���9ɜ33a�4�#
�h�ii~ݘI�M8d&��<@�~�aJ��6F�1���JY>e}	t��0�k�=P��)�񃃡�ۣ��4 f2>�8�#E���&�Tw˥̮��n(��4���`�=�����w���>�-�kM8��D9)wB��A��r�)���eVV	�;an����)�P,L̵�YQ�ՄQm��k"�ab�Qf���eb6U�u��B�gw�٩bbZhY�F�:C�J�ѩ�ҡA$i@�V	�ߪ�}s>%��g��?m$��t�Ѧ�K��k�������~�y]�i���Ŧ��S3v��$Fg�Lk� �7H�N�9�I��!.m���oy�^�lWp����^7.�/��eo���Y�y⡴\�Vxs~�����@侢>��������Fj�s�ne�M���c�&��no;��$ظ��)W\��qW�����ƅ�x���є&�ž�X�����/�$P��[Wr#�?���?)�YG��y��Om���4����:2��v��]�t<֘ȗYu�_���i�z�0��G�P0�H��`�: Z\�G��f��ą*5d������'�Sa	2w}�8uǏ;�l��e��ٳ��(��q����0d�!c׽�]��f�|��F�!fh��y��}�pBmC,%fKX�~�B�^b�0��-�K5�قQ�O�45ގ�9�MQ^�����Da�Je�SC(����>��E�\�zSdK=���yn��P�^x����.%ۇ�4dI���u>�F���d��P-��7�0�T\y�<�*L�7�0�u�s,yڳ�/��å8l�Z��p���������f���HR��n�6�������r}��p�C	�ꏏ��ٔ�>������g"�r85xk��ETI�Y?d��0� ��;F�JHz�a��~�<����i&�[i���ΚFRlw�.��2;�k����/8N���5��<?�^��N>�޾��2�ݦ,H@B�Ѷ���掮�C᠉���l��H�g�O�mݱ��e�	bF^qtόїԁ6d�"�; &�;��̫���N��L���;z�y�t,���
K��=�x� �9��ч&�A�B~V��o'd2�"3~������V7E��WP���(���E!K����.~�H1�x:����Vdz�0���)cpf���yt1!K��J�Z�����41�7Yx�����g3�v�s�O��$�48r(p��,�a�W(8�z�¬���<qs�҇��9��˯���it^��������b�%�DрQ$� �1��y d�����Сok��8��	
4՗7�ݎ�~i@���bF���̵����q�wgl�76�kn��i�1?ņ����CE�>.��7�ᘸ�`0i��6o�O��:�2P˚��v��v�j2|�l�R���|Ug{�]"%�0�/�P���3���gNy��Q��a����HU�iSI�A-\�����������/�z��vMh῍��ӡ���>��wJP��z�,�ώB��r�*v�t_H=(w�܇�=��C�O��cO����d�kOL���;:x���}L��e�ψ(A����1��$:Vǈ�z��G�Qop�s��:?}�	��\C�Ü�Cy9���^>�0���&�"	o�x��t�0� OMgpH)ø��]j8�7@�.4�k������n2�=]��q�Y������6K��c������[�tцf�]��c���3_��s�7Zxss9�j��&�>m>�Q�t��z��z̶�ٴТ:��oJh�k�j��-��v$�e�cRݛ㋃�N�ЛWkq�օm�\�ۄ�;c���g[��'t�,���n�=���A6�3ō=��1�Z9x,'Jsx1�P�oc��C[�f(�E�r��L��,�Dr�n��z��v64�1�w}$-^A�����ޏc�B����U����!�=��^��U����C\7���ρb�Q\�QXFZ��bv8�{�B(�!�|akc������6�����]�3�E=5N� Z;��#����r8���p���@��RK�O$j�(T�4Yewm����h@��v>~�Z����j&?[���d�^�!��W��;��7��	JөC��o�a�o��e�k�9�^���oF�_StsG�wύ��XVQ�k`h<�p�{�e+�߸}{o�,>>��-�|̟|�iʶ���cn
�2,&sAR48������i60��7݃g�P-�!��p�(�#�F}}$*����扭���q�Y+ۓ�{+�d�bD�;��!q�6��
"���sP!mR��G�+���K�)
h2��A�aD�	ӧ�Hl(f�x������^1wX��}�w��v��(������A���p�b���(�	�D0ܧ
��p�q��|����"o�3��4������2&��I�WQ���t͈�B�=Z�̙s1�UV���P���J��VCy���r�G��װK,��'��VV�A�;���C|��3�E��z�{�����B���t�j+c�"%�_���6`�0���	�����=j_:x�M�/��o=9��×��᠇���Q��sS�9�~4z��E\���T��e���j���<t����������L���"3��x�b�٪L��0�v��F�wC��!����Ot�#i�M�XBŎC�G� � A�v!�dn{qz:ş�C���*�L��a	��5�F0(\p8b�9����z�{��o�G�	�v6y������ܻ���}V�\]���l��[�����27MOSA����
�ػ,>��Q������8Q�@���B��"�ly?E���J����7��ƛ�
*a>��ߌ�� �5���w�BP�U�\r�D���t���Heo�w�x�艍A���T���Lg�:x�ʇ��x���8�M�0�7Pf��>y�5�/�K�Rm1���;��������ݚI�͇��w�A���p�5�v���і�ݲĨ��<ɳ�*`�5Y��U��U,�Tf�P��;b6mL�6N��"M�g�����M1�W.���ء"~���!���tX��!��!6`D�RXL%^8/.�}�>��t��|$/�c)����b@�\Pӿ3tsD��ϸl�,��GC��r{e��a�����Ǫ\�i���v������Ƌc�����}����t��,���׆���A��z�g�>�C���o�|�&,�#n$+����4uSs�\��]���Wj�X��l����/9�M�Zf݊2����ߔ�����Flg5��B�z#R�z�7���z��n>��{\58<S9�֌��U-�6�چY	0�� ��@��xh�^=������A!\#�C'�V�g~����h��k�PF���p�/w�=�+a���,���a�ד,�;���s\�[��.5!UA�?�s�*7�џE�r�!��K�!^8��`��Ƅ�Yc��;�Yzˎ�p��ܙ�S��8�;�7!e�.Y�S/��w�7f�orr��gњTg�1���ᆴ&�M8m#�i�m���M����Lo��s7}ﲒ�2��*'9s5e4V��eK��sxȵ�i���n�$2Yĉ"5����6l�z�b�Bwvq1n�$mؐG}�,����2L�2�]2���E�އ��A���[XjZ����Wlg(��T]*��������|��8SD�^~R�,)�h��y��&Ҵvn]�4Xc�����ؼ�^$�%N{��Ȋi�\�HZB����!�Q���h���>_�F�j�$?�3��D�P
���l�y���<~��h!R؈��|z��:i8�X�A={={��{_���	�����&a�u�����p��1�61���Æ�������$�a!Ex����V��v��ڝl8�Y-�.<HC��|l�;��
^�CH�Q�<���}6&��8�4}�C�e\*�hq}!�Iнb��Gc��S �h8d&��,!v4�!������V���U�,nu�I6.we����;�0�2nt���z��A�H�8j�
�1f��`�E��-����Xx�j��Y��I��l��Ϊtg��V�4Vi�C������ p"�S
(�ꦹة�Pˌ>q7!6��>���Q���7��u�����"�@����(ơ�g�wOj��0�4�ߛ.(��v��v>��3v�l��E�UVe$��=N����U�e�FU�]�urM�Зh��#WR&��cjlf�.���f�ho.�]�]��Ms��0����ޥ��e���l��B���./[��C֎�+u�Z��m�M�onJ��l�4�F:��8uV)d�$u�l�m�6!����Y���@��'n�&y�ج���-}!l�_�h�>��ک�E���O	q�a��K�3ut��#l��S�����,l�e�ш�1�D�[vG�_a��rUqۢ�|g�B�3��Q��tZ ߎ��7�,����o^�Wf]r��ˢ��0eltx�3"zuT4-&�A�Jm(W��0D��ܸqs�w�0r�۷;���%67N�{cY�/GD-C�C�|j�q�
��t�|YF���f�|�~,C�y�^\4o=F�YFbG*�U�����8QG��I3������k!8p+���;�)p�GH��X��c0,��ѣ]tZ�5㴫��m��	�����
�{�i���!p�z��D�ΰ�JMB9�PB��+�ش*��G���7����o�����iM�����6m�m�֦��!�����qj��!ޓR�!L)t� ��e#����) kP`�{��i��m���Y���r\T��5��$m�{Uq"l������:��p���]�)Ȓ%��ﵰ������),D�����!�Pq�pHMGl^��x��9}�W�����>��o�K��T(	�P��4�):�!:Nw�I/}�$_3_Cmi�J����o?��Qq�����3Je\��dd���ն��bj:f��RP�#A�ڮҨ�9[��Ƅ#,��3@(@�[@mB 6?��Ʀ||2˼�x�G�<ό��*Eg����!���K�$ga��ʆ����х2�C���z����.�$$�@7�6�{;�>����o
%i��tv��j]���s�o��[gf|<<d6�r���>ȠÝ<Y�A��s�����v�bAr��$#��4*=ߵ�RlȢ�@��r34E��Q��Q���>��^���?�e���*z(�9��e�z��}���$Q�0j�h��4�a��a6��by܉nܖ�TT���cC�21��#ո8���{W�z��i*��[IX��r{���bO�hjy�<k�l��v}�te��s
������f�|d�y>H1�� �1�B$S��"�����"!6+��|��n���M��d�r��>��?5��ﺯ��8����>>F�r�P�}���	��V���0�� #nq��܅BH9E��tHo��V����>�Ba	x��(!"M�#v^e�H;pf�]�P��L�'��Tj1�&�\o�#��V��3�k��ʐD��W��̍��DB�6��O�L��C�)�����	���X���j~��3�"��!�6jj��ٯ}����V��Uݸ=�2��Z'���&l�T���0g�!��Rׇϋ2�AZ���x����tl���`G�w�9��0i�&,%�O���*���m6[�C���$(�d@�����D��Q,z�F��vm/|Q��-R�A��0��{Z��{�����m�d:���wSkk���hN���Z�x����^�Ǜn�th�;=1����'o�w\}��9gafvx��oD���y�3G�/�YQ�8��~����_��W{��qr��}�!ȵ�#�==e�$�K����a�*�w�!��(��������rs���Z)�B��Zg�!>��2ϋC1�Pɟ:ac���|Xa�?���}����㉣	�D����1���w�7�;�t7L:|C�����ew�}��٨�YB>0x@7s�]�W��2d����τ[�E�/\�����a ��n�]�F�<^�f��8�����l�sd_ߩ��	x�@Q�����^��w?�@#u���z��	̪�)H���j#a:fѣ��IP �gi@0��cU)�:�s]�g3=���b�F������(HAM�e1��7�>'�Y]!�߶h���Ҁ�9�V�~�۬�^�͌�f��f���h�s{9f[|�3�`�`�A![��Z�eA~��ت.��@T�Ƅ
�����ruW�^��nAK�.;*=1��~�������T%\�wnꛪ������wVo��!�\f;����v��g��x����y��(_�
�X2(�{����(؄�]&̶�����OY��y?�O�A�6��3�m���^������n!�/�2�TS��Bٹ���a��O�G�xf��zg�Q��}�^�z%�@��X3�]�N#�C����ݺ:H��,�#A<1�����~��
4��4�6r󄅘}�F���_���S!i�]��}��b��P	� _��$sP|�`����kl}6Q�3X�-`��ѽ���7es������s9u�/��;��ώ}��!$wnU�p���7�@�iXY��-�>ȑ(?NW���0c�XHf��g��*���tB�:"��p���;
J�1Swi3W4�a=��dWzA��0�B+f����g���r���W�ұ�V٧Ղ;k#�`���;:`��aq�O�,ƅ�b�.қ�ta����^kL�:+u!-�+.&Q�ٙ�Po�-}ԥ����
)�a#W_�f'��R���lF�Rt���{d�yМ"�c���=yh����q�[in@^�ۙ�N�=
��m�<i���o�F�,X��l��ʃy��K�Þ7>_vs�~[	���t1״i����8W^�� �}�鮘KN�NYֶ�&b�;[�_V1'��9MS���Ņ[;l���ZU���*����{%�����iݦc��t�b�|�J㝺�qv����NUT�<�[kf6���:9^g\����V�!��έu6k���X�B\Iu��B�#`��s�_GZ��8�Qb8!d��;�[X��������ǋ4����9hW9�'7��)!�
��݂Qx�-��Q��P�*Tsi�	f!r���O�P�I��8�ï��fNt�Rٳ�r*�4Ȇ��,��}$]�78�|�Q�f�rz76q������[�f�2G��϶ElZռ�Ri�Ȓ���G������<�3�Ȳ4�����2$�.PN7�����(��?A̮n��(�l�I,8e�8GO��ZD��Sٙ6�ʭI���1tS�9���O`��(��+4=3J�g�l�EfGC�Zf,������?R]ǳ��}��@�D]PO�Gg�?G-�� �}�X�0@��������F4���7��)��te��aD�k�[ʪL��뉍��^�U�b�v7�e�����E|��t��2�J/�9{6���2�ν�ۓp��3�8���<mض��l���Us��d��4�-���S0�f8���:�p��<����H\�m�x�Bc���\pӛ�;<��ك��q׀��onQY|)l)@��j��#V$�=�}�Z<�;a��*�9շ����Kv�W���}�����[����բ+7-���hņ[�\�іۍ4R��I��p�t8�k�X`�eB�dئ���Qљn�y�5˄v�-YJCk�ڴ��ӂ}&��g�X}wk+ۮt��Ne���v�<���$�
�7�]a&�ٍ#�C���
WbK�O&4�ٔ�)Q��U-��]S�0�����uۖ]\�c��97/���7�#��$�6�ui8컆��9�\Id��X�Yn����v�i���[��x�	u�dܣǓ�k�X;b3�t{9��0�$�z��!�2"��ˏV��oRSK%#-���t�̩��CW\���%�3�F�А��B�3:1� �b�c�W���V1�z!x�$�u �4�x���Z78�����7g���B���s�����ň;u���õ�ώ��1h<s��d�p���6l��Oku���ȝa�Mof^�6|E���Y����e����I�un,t�f{]n�u!��\ri�k�\�ڭf������O#�̮+�lz÷�76Q\�v5�k]�&�Y���R�1]�H���Y�;<L����'ٽ˃%�b_7��5��X�Wl �vۊ��u��*I�
�ʓ]�vy3u����F/��m˺^�{ ���E�]�F�k5�b��N��k�5�ۤx���/&}nC��G=mz9����n�l���8�����q�F�n��,�B��,u6jf�q�oXBQ�0�d�s�쬢���k[7��nP㴻����yrF�my���|P��N��Y����Q�;b8�ɖ�nÓ�W#ƲB>�W�ĭ���x�n�+���m �:.�E.]][�6��~;4��E�.l�=R�/0�/�8�� ���q�U!�m��~�~wO�:u�r�>���lt�|��+�;+0E�ts��3�Y�v�����;�0{*�М��}204e�o۶����U
�'m����f�)��� d#k����[+��ZnNCP���)?��'��{v�n��8��/�~�Wߧ��6u��!�ņ�T��-w�~ΛՆ�9�|!˲���Z֌�~��,�'d�i��H�RH�^1;�;��8r���ǷD�^u�8��=ugѻ<�c͵�л�O`�St�\��M��$��9(	�I���t��8�t�ۃ(��w8�
�����q{u�B�z��p�S��Fݻ:@�n�)1׷>�p��X��T˓�X����v���y�q�7�����{s7=�^+Eyt�lv�\�!ۭ�� ���Cۍ����~w����a��(h.�,��Q-A�4Hi�v��TGl-��RJ&#L���a�I�� ��uRMm�R�2��uT�V���˴�
!^��Λd���U�oC�fA�w��!f����N��wR�}WGal�x���' ���$��i%��5�n�7�A���S��
v|~�1��a�}���,g8=N�i�9�G��$V�cGKx�w��^G� �7��6w�P�fDI����ف�0.v���a�dNB�՛0�r��{3�x���D3�#l��ob0}"�����4T&��Y(0E�g�ỻ����E(-���]�m�x(�cFأ��H��O_2�k��B!�`�4/Ѧ<g��GB�I�H@�.\�B��(�		��@H@]�&~r��P���|�+������վ�*�j���r�\ؾ6F|z�͘h����}[�t��Z��[������%��tu�^|�v��l1�1�����v��s	BU�*�"!��pi�a�*��|��)!8��{���"���o�vk���6�P��q�i�O�C�u�x�w��Dw���1�6�҉�a����	�X0�����_o�Rw#�mX�9�i���F5��'�j�ʩ�9	�.�+&_�䪿d�<5p3:�1B�w�dwV�?w�R"y<x=�G��" ���MѩF�+|�]dE}a/����]@ G1��(j�p���:�dO��4���`���^���V�f˭������t'�^���"G��X�0j"��=)��U���y��
	@�1`��  �7���(�8~_d��l�Z)C,$�^d���z%M4�"x�b�(L�m�,�>�,�������n�}�=,`� �}��6�+Ƕ0$Ĕ�%�V�a߈D3�����m���o�[�f�]�\:#�6��Y��l���� ��4����/��|��\���ƩM��b�M4�ܼř�hA�5�Z�&m�f���������p@s��l�ph����}��H��!j�e���+����Zi�؛<�}#�'61��V-4�@�k���gկ����49�O�"mBӒ9fF
g^�F�ۼ��J#~>��>����H�!�1����5[O�ݘ�{�:�7���׎ţ�Z_?x��\��u��G���C��G���
��{��q!�������=dVύ|�r���cI���|w�wFwF�L�ޭ�:B�Kf��)�kUs��UK�驠G��xv��'�� ���]����+�@������Ӎ."�a���C}����ad+��;æ{�A�[+_rk�=vU(U�����>5��x��w�����WK��pR�������h��t ]��i(n�yt@�-`�X������{�.zϏ.���=��Ώ���Fp�D2�J5��@@d��zX�,!Aua�J�N�,���7�y#���-?��p��0���e E����9�g:����5C�Uv��+c5�nm[�"�8ց�.�.hc5��@��h��AEĈ�D/����8�A���\x1GH�D�'���I�����k�ctn�rn�j:5�VH�n>R�띶|��ڇ�X�$M�XC£����
q($���ӌ�y�щp/���j�"���gك��4B��@mH��B����s�OJP���]�K%4�Q��KC)d,�]��a� �����g}�~���S;N���dV��<2}ߞF���4� mW�/JP��m�BD����1�6�E�X��k��|�g:;�d��_s�xP�VΖn�Wāc7�"x�J�~"^H�`���u��D,��q�Fky�s�s:�>��}�<.���//���^�$��fE��j6=�=>	�D�jE��J����!���o��X|�o�I�%	�Y[�Փ�
�!}�k0�/��4z��>hp١���Rk߿����I����f�UD�[;8��Y���6θڐ�;Sm+�ˢ~�'�<}d��k�v��(f�nR�å#ƠɅC��4Uwm��M��<�ȱ0g6 HЇ7�FG��!L��@���á�层�^�"E"L̸E<�>ǰ�bF�M8檮�c�Y�>�K��a�a��C�������}���:��(K�nE��/��gO�����-������P��v?�K�Xa�0=��=ӻ:���F��1�Mpwg�q���&v��8�Bz�@B����;�S�R��aƶ��`��
�\���0�H|�(�&�i��	���?� r��d%�f3	K�@���zg��_(�M�F�3�la������K����B<���&�XB��E F׷8P��o�,��X��H�I?y+M�E�̱k�2(T ��walܬ�QX7E�w�WBd¶ZK�gυY�I�U&�ІG ����LhGE��:�\�^��iy6Jg�iQ��\'c9�:��F^˪�1pɬ�2�+v�K�M�p���V���i���\bE�m�O`H8�s��^lY�(=���-r/8Y�w&m�f�{7�]�]κ�r���]s{�x�ݹ��km����K�#�Y��*��ݣ="k9e6pb���O&�]b9{t�;Q��k����D��7�˳&:�3����^~�������'3��tN�8�>��<��;hX����'����h�X�.�ِi�M���u�|3���H{W�5pi6�1c���HK�����h��4I��H$�H䏲�T!Һb!�_7r�C3��Y���G+ݑ�Wm�J&YW�P�"��s�7�����wf&6�������!"�ū��P�}J�p|��,��sr��������%ZwRX7���<�׌��}DXhV�"���C��k=������<Q�D#(�OR4�����
8����}��L7��b�<:�!6���`*$�'����}��D&ņ�UU珆r�|q���j��LX�������=!�̺�K6_����<Ć�����rb��"�{�#�cچ8L�=�����Cj��"Bfo�ճ_oFa���I �@����������vF�ا�����t&øW��س�/nζ�%���Oz��ަ��l�ƶ����Pr�ʬ����e�6�Ρ2��2���������O���\+�}8;�l4K���<���ޭ��'��:`Z �P�o�1���UD�eP=9�P���>�ܗ�OT��Pӏmv� ڝ��g�5�S:��W@ҬQQWBڦ��!�9�G���iK���.��a_/��kCsa�%T!(r�ï_���)Ө��܅��ڜLh�Xa+�><%	���	��1Uu�,S{�Yǘ8`�Z�M��M)+.�0��_�6:G�w���0[�X,��o��g����c5��TN�h9tkm�(�g���� ��6�ۊCޠ��֊��b�6����,9^�պ�4�M	(���7
Y{� ���fn�e���o�_��x���������$�(�p�~oD,65�E[m�YA�+��L�6[K��Cue܊ʌ��L�4�+�b�3t�B�e�\Wm4�6t��	���.̥�TO�����d��7�����.�=����$��(���LmY���/6|2�tK~<B�٪
c�s���(���N8[-��O& ���o�߾�F�C��w���P�[>AE||C�0��_G�5�D&���B�4��7>z&�3Ύ�j7v�T�J��9�!������ >t��ψwvQ�Ntp���?#^[�ll6�lQ���Z�Ad��$nM��>~�x�@9(2L�G8m"n�3`l.ۀ�
���M8�"��ܷo8��LЭ���UgW+���}�蓮gk�f����ck����aÚ;4Q��G ��P�ke(sː0���"M4�B�}�}�Gu_G�:#F;0p�|p�x��O����Pϳ����_-{��ЉP��M�c�n�����j��IZ։��ڀDn�D�!�-�B`!���2���|uxD�I�l��x>��Ej���7e�q�*԰m0��6�aϧ��_�?��Jm��mr7b��:S=�խ�xAȻ6��`��8/�������߽�|����6���KS��"�����W��]>�^}��d!��<Q�����]W><`��������(��x�/�C�t�~��Se��<8��ώ�[!�4C��W���<�W�V��M�E���C���f|Cej���_	)X�|OQ�<H���Ki#���>*/�4B�����|8U�ۆZ[���]���t��<ADe}!���D��*�t8A)�:�C��ē8f}��u����Q�D� ���?h�A	4�sXC��q����m#��o�u��.Q�$�]�ä�}�ݤ&��1b�\���nM�roFE70'GiY�Z�����AQ	�w��o�X�c��]��kZ��ߗL��fk�x����ݧi�Qې��U�G�t�fr̆�3� �/"�BI��|r���'�ᅔ2g^�9�ٛ`��t����n��m�ccc7��@�x������#Im�1��A�ʾa,U���mp�l��!��Jcm�[O���}v[l�N�uD;Ӄ8j�~�::3HC|w����q����l��}ާ/��s�0�r��\�咎a	��:d����������c[��|̉�4k�/�+=�S�P��	��{�.�QvX�`���uc>޽�=Q��X4_����5�p	D�s0��P����֏��j-$`(��� azj�;�0n!T0PA�	|�D������S*��Rr��r��B-eP����� xe���<Mt����>!�Ӧ��߲e���nB ��:7�_�P��85,���}Q���HX��Ұ{���{�3�v�|0`8��1"B "Bᾞ0�AE��6�iT��ދ$<2Sp2�����%\�2��>�@Ad7DLi�{f�D'ܺ����Z�C������#R(b�JT#dӵ��]a�[��X�)�m�B�1jh|�n��H�O[�<iܣ�F�r���O�ܜL�N.{T�q0��`l�6e�b����4l��ƶ3�j��g�Yrx���<=��/\��ٽh۳�ϕ�ktn*��8�zs۷	k�ލ�-u�{6T�k<q���	��*q��9\��7gmm�.��2�l�b���R.K+��IJ53�2�Yܭ�F��5&i�'�����զ4�\���;�O[��vdI�{tɱ��gz�<��#t��ŕ���!$4k��,qt�|o�Ѡ�C0 ��@z�Vx�r9!S/�`�c������I�,+*8l
$��P��@_`ձ��y�&B��z0�t�jn�x�1%	GK�F�=hp��zB���'����e�An.�.\n�h��U&W��[K�0bbcq6Q����:Ye}y���<9�3zoj���_O���1&p�Q�g~7%��&�p	pa!@��[�@��C5����}��٬9j�Ms8��xv:�"��hЀ�A��X?�g~į�)�څ"b�X��6�>���`�<���B�����<l�A�!�p�6�t��B�m�`���٘|T+g',�M��lhh���{�FO��g�R_+�sX�Qu�lq� ��o����wS%dy�G��mY�~�Z�p��I�@�K!��P���[,�WD�o�",!C3����ڢ����-}���5 lmD��G����0��."���hB}�p���Ǎ�E�$��(�]�n�<��r�题��Dc..T�j�g�N�l�7��nb\���b���xM׷'}�����8�%���{�K�B4���tDh��L@j�eD��n`���C��V��}��@���Z�ve�����$/�����a��Se�r��Ot�o��=~��c�׹DeLZ(�w$P��*��f8p�*����~��$��C~�<�Qo(s�L�	6L} �`����t���5 �<4��q+gFg��������/�f@�UE�� U姡lW,�����=w�7Ӝ�;��ͽ������K������+��69bw"�H0����-�A4$�M�\f�NO\A]��{f3[�k�����e�H���ݙ5� *D�	2�暴~�xq�]����x�@�b���<5��s�|�ʳ��e��yt���ɾ��(�q��	�����h2��J]���64!@b�����<<�u����gV�@<0Ƽ����w]ss�л�8:��^�_{�d{�Ћ4�(!8g��y_t�ꪸ9y�9�j`��p��NN�?����	>��`[��G�L˵>�xzg�ě���v���gЧD��h=̟p�c#gd^=f�I���3������OG����s��:܀���s˵����^V�-�:z ��ι����8b�K��(J�}I$�}hKu9�X�{�7H�����.y`U���ڬO6��Ҳ=�Z~�#Tr�6�&zo+W�B�sS�>[����P�r�ά�z8�D��]L���nV$�:��M��[B��{^�?+��W5��@�Zw7�6�=�tg�j�1�bU��o�n#f�7rΧ�yU��9���
9�$y�7���kvf��9��"��x�WD���f�E%t�v`�w��ք�ˇlp���r���uA�S1�>���p�6s���f��=B*$#�t����.��M���(�V�٪w3ܠ����՜MIh]�ˑA"*����#/�������c{
qz0�}O^ӿ��r���
�xOQ�3�o�_9��Cv�	��8��6��"f�e�Ƀ.�튧�Yӧ/�.�LE���z#����|�!^�8��W;/4t���^�yq{=s�c�]�Q�=-���^���$��q{݁��.�%a�sy���j����s��`�z���εIdgN��1�b�^v<UU�ӓ��<�$��h�I�o�jq��ZҠw#a�����K#Lk�)�3R+n�_]�1p휭�� ��JS��y����I\�r�Ÿe��B��=���|8�Y5"��ت�d�b'���l�ݵQb�����f�<�u������Pț��3��\�b(N���UQ�	AĐ8j�5/������Ol�����6TGG3E'-=�m���Og.��hu�Ze��ʞά��������ځ�Ӵzˎ,�']�/���z�;��R&"8�8Z���R�h-U������;/(,��R�U�|���NC�I�F��O��������TDD6
���L��m�ހ�� @����%�ؾ�B�>T}C�w���NHT#(��-6BP���� �Ec�Q��Dvv<Q?��~��~O<z<����L�����&s�r�r��^'>ݼrIC0��(x�0��#g��R�<I���U����[�wg&����d+��V0��t��	�ƌ�a�al2�V9
�7���6v�sUc���f�1|n�X���Ɋy��|���!��w�`�M�`�L�]0��ۉ�%�W%�1���{8�6 OY'�L�(d�Ѿl�d;�#|]��wZ����N٘\˶IM�'�����?oǮ߇ט��������lp���w�����J��BDI���^�IAq ���G�i�5G��1��^����f��}�i�������ad�����UU3�yF��G*�m�MM�o<�<�hTj��kz⫖\�8�D��<���Zw���Km�݇Ua۲��	lx�����#r2�gH%����>�ߏs5�h�<�M�I(�M��7O�!F��!ax��*/ـ�}ͱ��I��L�0����f�ڇ�Z�@�?C��/����ڻV9�fz�݃��t��8�n#n���eܤ	/i'��i�Z���J8HE���?�\(�����nK���ͦ�i6�,�8Fs�ײ����nz�2?��'�/�1�1WfZmH[������UI��\��n�+*��rof�'��_�6�Q����O�״�k�j�N+.���A	Cq�P�d{ܣ��:6A.��gzm�*��z9���v|Wïo��_��yNUeU:˂I��g�W�ì=��ڹ�F�C\\�ݢvg��YA����*�=G�&��;�<A�4��e��LGI�O���w�!!�i��i�lq�Ƞ�^��D�'"?�"�����ũ����	��B�!{@�\�G�4}�lď��5wo��6�|�\�����I=CCl��P�5�U.�[�0��ы��\���/�){ړ�c�Uh�;�Or�v]��XW��G�i�3�i��d�gIuх��5�z���> �&9|��F�:���ebZa�5�d������f�.1˘��{*��\^+zm�m�D�ID:�Z��5��F��u9d��^�s��u<���]N�[y��J�\+���۶�-�،�9W���a���;�:��eM�<�Ļ*���X3�n�vy�i�mt�{C)�\u��n����%��b(����Qm�差l0Uy����R߰~W#8�M&�i6K	Ԗ�W-Jm�����k'n���l%�i�!v}>��[��Ҋje8�	�C�!�$!+~�w�!��"������'O�9;�����A�����ʟB�&�L�d�w�r
��z�*�̮mԌ�PH ���HY���C�΀������k��c'|Yk�c�ޚ}�t�l|f�\P�շ6��5�zU���+JMo�m�^5�<�8P��7�}���>#�wް��i�!�� pR�*��X27���!>���
���{�{
Ɂ��p�T��@c<{�|D�	��i;jU����N��f�P�ԸSd��ԇL|(���p����BlQ|/
�HI��wew��~���w� �r�,�I��3�U�u�ɓ����=���ce�N�9���OϿ9J�lɘ/�G�)�?�����v�EA�ޒX���|�T(��rf8X_h=ȡHG�*���+���)�KpX%�51�N���h���B��P�jS�&F�3���U�T3�٢���F��'V����}�
�Q#4f�x�[�׌I�(�5��tG)qf�,䡓��\߇��i�ha��=E�&g�F�p�b��
�����{2;��=l�%\pd�3*ȃ�a\��3[|_~5��rY3�\��5�&>�#�3�_,�6��(8%&�YM+��>�?b�z$xF�_&���h�A�l�L<c�ǹ�(ǹ��V��aOl��氭w��٤u����;j&}���J��%\���a}���m|4E�f�p���'�_��E`uN�C6��S�7�Ydr��$�|�pjB�;X�5ٷa��J���N�lc���wt�6�?{w*��$RN.�QC��}����b>��H7�<*��C��ˢ�0�n�PP���-���$��-B*���~|<~.f2��D���;�0N%����v��}�(��%h�k��F��e�u�*G��E���;� �v����P���ӍG��o�t�/�/�< �6���P������G\�K���vd#�9VeS����B���G���X�>������Go��M����x��c��L��?(Y0!��������988b���{�\d%=��?8��	_\�j^��s�uF��0lH�	�:=��w�km�)IR��Uu$��)=�E	BҪ$%���Bs~��Ãv-�2/G�^�rNe_��{m�.�����J�[ԭ�V{U�����K���6�bri�[�غ�?�Ϸ������˫r�eG˦���Ø=�gF�E�||fu��{~�#~`*�(��d��OГ�,�($ըF֊>		�6�?\�q }A�d�X�)е�<22pxpbFTϬ�����z3�H�����*�x�ɫ�RP�|Y�a2�Zȃ���戏�$H������$`a���&�#�_��M� �D4l�|4<���[���hH^Q�Аa��l �H�%�!�'�r
*�'�4yO����|H"�����O��Z�Yg�x��+�|����d~x�S*OW�#��4�"\0�Pq��k�tM��]�gV�<�1����D�I$H$�*���Y�J�W^\uS@ރ�Ƕ��sE����A���@�z*�}�,3,y��ɂl!�C�
�i25����<���.\������w"[�A72A�2[%�d�<�[���XFn�8�[9&&�Ŗ��S;��z��K�8E@�hWH��]�	o��P�\1���K�n�Y�}��q*B��r�.+)[e~�xy�s�>zy^���Ö�h��̀��� ލ����(z��|(�rc�l�!3���C��)�(B%�}�#�|G��f��]݃$�%}~��&<�C����愄�|M���yBi�S&N�
e��O=��P5D��.0)��!��C cV����r*�<�R�����5CM���4^�o�/= �_����@($��E"�"pк����Eq�|���7�@�"SYd��	�#w� :�!؈w�c�A���K+�їN�U^x��E�F�1�,O8�����xnf�;09��CH��4��a��l�Mp���I�D�ӫi�裍Z�4ghWq�*'��{b��=5�I�a��V��b������U,��mk�݀��)m�٭�f[bU�a���hJ:�XQΎ�i�����y�|̭����c�Ux��Զ����hړV.̦Q�3���Kp���V�\UZQ�s�cK�6lN�O*�lt��<u��B&y۫��8��W�K��]�oMoؽ��ą�Nv|<��$�':�F=��(�r:�ĥY�tz���n7S�.9b�a����w�a� ��	b`�B���hj�������s��)�UX1o\(QNU[���7d7Ի��I;i�>��MTՎ�I�_g���9ރP�	�"�W�ݽގB�oF!8P�8e6�	[�/�&�8�ឋ��G��������Pi&����P�M�B�q�Z�(�i�C�F{;��FL���ӫ�6Qn����ٳ`�����~g�H�ǸdO����K`����	���C�0�AȱB␐�팁q�w������	ʱ��tg���b�sK�R�K����	�=�Ӷn�;�J��t� �#��LA�c%!Cc��7��E,*H܁�f�P�<��2�U�{��9����U�N�N��_����/�?��Eyv�p�����O[�N��B����GƋ�^ȓ$0�4�%��}�{��"�N`Qś �:�?�6]��u�i�z���׵�&_۰��X�R�+��7u�٦�!�UG� ��2~c�Q灝�R�
�N{�L���ː���Ɉ���i��(=�J�
>�Y0!�/����z�\�u��P</����'�A����z-(m@M������cӌh�K|a�D�Z���\>�0b�%ȓc��HCC�;�?���`B"�}���U>�a�0S�)3�������_B�R=S���P��0	'��~�������/�bf%-�i.��W6��t����2�4r�J�#]\�DnƋrtF��1�����m�_Wc��:4�/�0n�r���Y�}�|��7f�I�q�����������K)6T�8}�b8N�O�b�OC�$sb����p��_���m�WK���QA�Yj%8
 ��i�q�{5��՛i�7[>�K\�m����m1@�	1��g>~��x����9�C�L��)8�0�!���d,(@�WFG8"5u�.�LW7��'�ݺ��HH%�~݉\����F����ON��GZL�B��E
r`O�S���-�J;f������#ȼ���|$C��Ϗ�<�|Y�@��Lf�"p�5p����Y�P�^)f�K��Cdf��!�����3 Ä���^���0�������#��
�~+4��N#C���$�/�ϻ�t��s�>k�������Vɖ��'S#`颣����4�]GI�,�we��o~]=YBM�>3(9��5��<�B�p��k��}Q��.��I0co�&�4;�L���i6ʏ��?\��A
�7ͺg�$Ɔ<�}�`1a=U�|/��d��mK>�H$}��[�.)��|Q�� ���������=rR�#V0C��b=�.`HB�>6u�>u$�)�<�
(A� ��} �a���ۙ&�=��Q&���l|록Ѱ�.���'Ff��x~��'Qus���OgF˨P�G�02M�̀˼��s�e�ܑ��ٻ�w���B�p��7�m�U�{�@䈠��6�\A,��nAp�HT��wBCSm�oC����� ����ppC��ʹ�+��\C#��0���ܱ��A6���	��vn#����\�[f��Xw}�u�,�y.2a/����M+Ў
���<>:�K54Ϛ��3����W!ӆ�z�|����%�4�vXz=�|?�߱!.;Uz�I���с��4:P�h��&�<3����p��!��y�XI��H�p9�GtV�f/!PXf0p#��������I-��i�l&�hT<����.�����ʿGڏp������v��1]�tW�kk^��H[4}���p��&���)< ��b�1w���ܶ�����<�(ib����xn
��3�z������[�H���ႬT�t�4 *�J�Ԩ�/�KfطЧ�=����L�%���8>��N��6珷|Z1L��>�����i���#Z��{��s��z��{������	�z����W���$��({�H�λ���^�{T�4��0�Ӡ�U��ϥ���s4C�:Q�̰?��W���r��Fw5��t�y�9�u$��ٍ���/�]��w��F��g�5�ϵ�����d2Lv�?�Ż	=�d�<j�6��"X u`�o^H�P�6nb������������
�f0n2k�A
���eN&w�9��{;	|��y;4���Uj�fw�ia���͍S�q���D-sQ���!]]��ɉ/�E����{�z:0��ъIa�2�eP����p���]�ԏ��<�E>��8w(�`��������-��sX��f>tu���F��k�emR24����J;��ݕ���zV�IŹ�7P.)����ktMC{ܢ�am8����c ��^j�f��o����̍��Rg���g��w��,Ɠܧߴ3G�~q���W�ݺ&W1��^Q{�LY&\�B�nl ƹ罣��fg�Gc;����O����e듎9��"��Or�W#����{��7L�:����R&pNv�O�%�e�QQ$@���b��������IB吺�R��srU�n��������/���k�b�j��'bH�B��;p���Z����r�l��G#���#�K����wn�܍ZT4���"�[Os�ػW{\��xYð��\I$�n[�#UݴV�u	D�6�U���q]�[iY����Wr(�`��$��fq�d���ۇ"��˷;-�qptd�Np煣r�w`�룎rv�^�0x�q�帍yz6M�;������/Xޱ�k=k��G/X9u�S��uۦ�u[���iʱtYL@��6��y�5�u�gK��S6jT�;cWC��X�!�N��t��`Mۧ�n��玸��ʷ-�V+z(L�w=,��g�f]�;F�n{��o<ǧ<8ħu3ȍl<]�v�ջmۛ���ܽ-��^�v;���eݫ����M�:୞�)�E��v�%vsk)�d�hM����2���݄y����vq���;DI�.����h�:��%]L��8�N�͎�4d��v�f0
v�m^�����62�6Ɣ�C2�]h��kyz�q3��M�]M�m������l��"9C{�嫣q��tM�S�ArxZ��ۄ	]4Z<l1U�-���n��[��nz8��y�3��e���跫�����/l�q �F9�6S�On(Z�ۮf�ua���lֳ�uv6-Kr�v*ۦ貗�c0̓��jB�=e�od�$��v���do1���� k��M�Ib��i0��ҵq���"���;v��н��v�v�}T�`�f����\��kNA�j��s=�*��E�(�{���q�p_dWҕ�ڒg��m�m$H��ю�O]����ةc�\X7F{.ф=�Ÿ���vc��[S#He�pk��U�K1He��
�j:Q"��6.G�������Qv^��ַ�on9&�����x\D`ѷ�,*`�y�-֖�7V��l͌�fqR+׋��KD��nL7l`����̹�gB�6]ðcu�T�<\9M��Xz�12��:Әٞ�Z&+�ge�v��R��U�K��`�����w�.��Bg9��Jt��s���[����]�c�3�L��Y��^׮Ů.�]�K�v\�Ϧ�[q��!
�n9��Q�\mLw%�LF��[�n��a�Mi잏�˖�ƅ�pϓh��7P�foD��}�y7�b�t������S�'f�>����*{B�74�uY`�����b�mK
��jb���if����^�LM���`��{�Q {L�#4���쌧,�_K��n��6��bц'Fm�ůN$���s��W��vZʁU�LNq�;&b�[s�ZuF�ɫif��]��[&�򁹽�+h���]nu2���\�]*Zm��Y��������;;`L�5dugt���[�N��j�dx�n��=�����gH�s���h�v�uG+DV��0���#E��T�:S�:�\5�d�tͳU]�:���&1q4����`x�&�ukW�N{��ATt�ױk.��Z�\v��>�H��BQn��igXA�-cn����ƛ� t�-��%G3rK���~�ٱ2�a��_�~��w<������Mk�v��a��{<����7b�<�ڷ8q������'�����F���燳��p����|��0�24�C��Swn׷\5p3HS0*3����P rP��X�?L-}[�g�;�<wFY}F|_�h��pEU��1]YP8@�/��AR$�@Td�ߌ#�B�N��[����+�nwb���HS�:�`��HV+��1�7��͕UR�Ie�R�=���G�I���瞎>�l�EUB�>�8p�؀�4�C�P�u�
�O�s{bD48���ق�a@C�*(��}�|q�Ct�G������/X�nȁ�ހ��+��H�,b��.���޴�h8E���MED�C��ġ�6pq�F$�Ć	U��9���	�f 6� B��ȑa������06�L}�ɴ��Gd7���{���I���X�+~��}D��i٩D�a_Nދ�tz��i��(לa�Jk�>�p�$a%0�ӿ�3L��k���1���0t��gfpیN0�ܴԬ�Qy|�9a)\��99�In𣘲D�F;GP��G�7���>������F{�$%�<z�#�F����GT0��G
h�B�����ޠ��'�<���g�KQ�����Dz4����R�nD��(�I��|�<{v˷.����*�G���=^��[��W�Ǽ���ᤱdx?;�t1�,9]�J'�+��`�1DBE��Tq�Z(Z0w��>�0�_���vt�����9����|T��ݔ��C$6�����D�F�ebF�3N7Y֞�-�c�.�����ZF����זa\I���7>�?����N�ؘ���9�~�~���*߆���n7XX#�h��,PxxI?�dO#�ʐ���Bu�`�gx$2�z�beG�������C�\T8Ͻ��|�q����3�3����Y�
������aQ��禎�����w���|5]��Yi4�8K_������qG־Iu,��J�8ZbZ�Ul��Eb4$�UG��Y�����S�C��w�����fX��������t�H���&R׏�:"��y����ـ� �Fod��-�F������㘊	/�B
¯�G�W��#`ؔ��P����8E0�"���ׯ9I���b�M��F+��΢�p��){��$n	��?S�6;7�ǲEm��nPTB1�Hm�
�l�LE���*W�>��Nݫ����1�~��]q���֯��������I?|��������H90s5'/�%H��	�A����M��Bxo�!�H���Y��;�K"��7����:k�WMV#x��_H��Cv�e�T8��0tg���o4� ��f<�M���E9~=l?��=�E��� �|���� ���BD����ހL(F>�ہhwa)8c�xx:��{�� �qo�n�uNꝪ�Ƣm���a����ï��ӄ���"�������Ӆ� ���ǆ���w4j�~&u������	�������.����4�^�c&�����_�+��jΙ��������U�%ݎ]6�>F��lb ��W�4��vdD�����w#�/�(��"!!�9~��[��=��(�p��$�8ɍ�e�;6��	�J
�t��A7D��D�Si#��%��P�.A�sV��0��M��_GG��v��p_S�6G�(X�Fjн�)QI�-�p��H���8{�7���P2ׇ���	��T��	j^`!ЂAooH�R��o��n�$�$�hʎ�Y��z��v8k�bb���A���l^����^���V��}흐������[b� P��9�d&��������mD��@��44� rJ��`[��b�z<� t���	�p0�!8!G�~�����gŮ�N��_�/��يx/��V?��5�����Ɔ��+�����y��,�9�g�����~p���llgH�;�]��O>�׫oY7�Y���6-iDw\���*��&�Y��?�"��$�Y�'(�j��D$�o�#[h�qj�(�i㞌n\�\^eキI����c%�����g��wn٩�v|Żuێ���v�j�s뱋X@�o �l{nf�nS���96���ìm��N�:�R���9�X��=F�K���>�5�綶-��xɈG$[Z�7�,j+��X��{=�9�u�Y��h��<=M�W�����2.]L3�
bLAjk�"�"2}��<�~��Wb7x��ب��^��>����l�
ck+,�宗W\�H�,1�9��1I
�D��8�p(��g�8N�h1!Uwn���۲,��k�<D�<u��g,��P���&g޲��<�����nS�6[r@�Ѳ����?�����B#R�@��E�]�1�BdxHOE<��\�F$|�a1?Xgފ���'	�l8��!�+�<$!����B�W���TQU��)����������z��g^;�M�;�:eV��r��K��٢��}�1��jL���X<v��ʶ�CDj����b�M�0sǋ].����|F`g`��8�0�G���!	n!������	��(EVv���|C�}���8K�	��(��6�S�O5���{1S�25��`���jV�F��Rj��:�9�f �D�E���w�fi\�8��%@�	[�� ��8]�PHw���Ҳ.�cc��f���?�N)�����n��8��c�wc�|w��NX�<;oS���`N���� f�q<.���U�N.#��R{���G\R�tlZR��EI���S��`l��w�/Y���fSj���������!`�<�e�-�0�m��t+�ާ���d,lI�c#w�t���!��|{cLm�����2���$*��9����^�^����*�)<Pc���_`��N�",&�f��};n�H��
B8��*�e����D���x�H�d��7��#����6߯�tHU���^�!-�ol�g�G�ȡK�+y�{����b��
$���[-��q����S�H'C���n���mѳ�S��+��-�P���0�_1�/޿�!"芽 �F�w�o�e�H!0E�Ho����8i�Ra�LVXo	�\}
`������P�w�5�4H_�cC}룟U6Ϥ{:>T�}��겥P�U۔QGa��D��=����`{L�Sᕪ���0�dC���i� �Th�6�g4������Yϵ�he.�=�
�WLI*��գ�a�+B��� ����LtF�_�+����گ�R�F�G��@P��!���2ۯ�y�R<߄1Ä���?T�/�>�+/�Ex@���� ���^��8�W��<Q���Fo6G�C]	���Οz0Sf"0�L$)�˯��Ov�*H����m`���py��;�0��Q��S���������Ʊ�8�k��jgjj�k�DKZ��M	7c�zh�i���]������=C��  �m�w��M�`����U!G�Ώ�=���>���Cc`��!O���Ʌq$R�A!X�P~��	:��]ͷ"���x\|��Ϗ�>{\�)wCd�I$���~zFs��}�z���E�~��E#��ID����~����/¯���W^�t'PlFc�B�}q:Al"���"��z��x���Q���"D֋�-
Ls���@�=vP>nGl{��?d.#���z�G)����f�����՝�f��}�!J��Ӳ�yF㙑6�f���G��"w�4F%��l,� ��o���!座z�K���Z1�+]�6*5�(��E}Q�8__�C-p�۝E��:tf�m����]�ʝ�����j=�V�I����5�[A��ơ��`}�ȡ[!�H/�Fwy��K#�gvЏB�Y�9S)�N@�r��w`�!	�*f�|>&<c��'>n�o����lm�496����1��׎�|BB)���#V�	�|\(����`߁�����	��*�!_Aĕ��JP��8w�o����Jb@��2�ꢏ|�ΆeꜮv��ͧbC4��!,�7�~�����<L$/o���fì������?C�KT@�Ի
{��C�bZ(m!�y�!�����6}�g��h�
�Љ�26�7�^k�p����I�9)�S\c�}��c�q�����CJ(��Ҧn�j��i�^"�tGs+Q�������i���8Ww!N�ed�ES$n;�qz:,��5؎-%m ���I�hS�R���F����<�]�p���ڣ�s9[e6�⍸c�˱<�f�Xs�^�����ml�y�κ�X�M�x$Ѵ�s���v��sF��^�왞
�*[����vŷo!�!`L� ��ZÑU'B�k�k3\�[eZ�Q����b�vf��-4�df�-0ԃ�]��i�ϕ�~��CYJ�*;��!h�p��mf��Ϟ�w^^�"���6�KPbrl��S�ٿ_��):�Lӏ�!��GiH�4g�N �k|��G�/f2j:y_*�잮C[���mAq�	�	@�dhfb�>j2��gQ�4X}^	��i+��B��]`=r��p��$��z���`�m�	�`������ S�btཱི���y��_�2=�L�.s_��2	z�$b�Q

f"7��[�T��ý_U��H�z�$|����_R���B� .#2�;��B�1�!�=c���䚑G���({с7~G�i�1�	t�<'�{�P���6,ja��zO`D�%MGn9f���0nF̖�ae�,�cIۄ ��Ha��#毘��[n5���}x;6�7޳�����K]2od�?�	a���AW��=��(%&�8E+�P�R7�M3䨡���Ȃ�� ��d>^į��.i�ص�9�f�IGgJ�g	C�nH����Y�-K���3+��"�pT\�u�V��{#Y��,ٻ�}cs�ֈy},p����"
���}����ކq���5�[j��/��_n����Jlr�e0�,!2���G�z�.���|ы��h�2�w�u �I�	�m����ޮ��x�K�3w���h�[�K���'5���	�}�6-�Z�K��C����~��G�=��A
DG��Y�v|F�0F�]`��z�"k��z�o�P�Au�bc[M���cjJa$Ky�g�Wki^ֵ����P�iZVVBᑧ$LD�������	��儃�3<���H�H�᣽�	��T9�XI��&	��;v
�|9/�mF["t{$PeD����I�=M����*�Og���u:"������%Ȝb"L�ɡÄ��(O�6�r	�(_�/��R�������uRB%�j�}"��ے��%K�n��-������*[�ְ��ٗ��}�.{y��y���Q%�Ax31�{�;�T7��#h$f�U�^yXI&R�sV�C�A��Wn�:����Do�:N�G��ʽ�XD�\�l�F�
��N��E���x˞{��cH�lǡI";��sFp􀿰R%�����ﶎlW>�vep:��h�f��ڋ���|��J��� ��7I��{+�����ڨ�cr����:Iջ�K0�g��_G�(��Ʀ�����#5e.�[�(Ɗ�)7-L���Jv]�&lR�#F¸ˣ��̮��p��H�Y2���N+�"�d�g��j6g]��˛	���0���c���M(X��b�F\�y�Tt���(&����We�r��W}J�VC��}�;wI_J �]�v�_P��5h���.��S�� ���-�|w���yY�a�\����MMcG���ԥ��׶�ŇH�$	g��0�5fo�D㑨�D�rcT���j�\w>6~� I8jQ���Rs)S��n̺�%�e��c�8U�}m�<�LD��;a\Fqǆ��ny�j�=|�Ft�u�����"�"v�n�ӄ�.���t�HjNU؞��z8MDD����:Z�O+G-,�� �Q��J����t(\TW@�(�VLKH���t�qY��Y�1ToHZ_N^<�r�����F�H��q��ƈ�zn>�t�|��N�k\��Tԟ�5"�"��E �0�fZ$�KˡwB����:�a�B>#29�v�g_������b�7��5x��PV�+w^;xz�6�ɠѼ�o70��$�٧7*��D̪՛���3#<�n-pǕ�C�����h�&wL�L!�.��'�<��g���ܝ�Q��<�^�d��a�����mi�w�&��f�;
ܼ�g�5L}�+�:4�������F�)U�T��r�X���%�oe��p26�[�zK��73�2��e����o�ý?_G_�Np!7=^֊͙�{|<ETg�� !\2��<�Yb��Q~lM�x,?	�~x����((�O�h9��T=l�{��/�����E
C��Ȱr)�P~#=链�/�Ǳd�K6ikk���nn����q34�8������(@Jq�?a�wѮ�,L��(��g��� ��އ�ts�C�E�a	�\7���C�xP�3������J�#n��'���Gx����1����ۣҨ�*is>��P��RE�«�� ��Mg�B#t�r���M
���E�
)@	0���><p�鲎o���~;�p�D-͡w��r8�&+;K�ـ[p�H�A�^N��򩐦(��B��TCʍ<7��}�"	p�KR�6C"�!*_2	�"e��Oү�=�`��.���9#4��!ko$ވ;7�B)N�*3#���Z��R�?+`��IŖNؓ���:��}���x$9`�� ��\����v��IV��U��1ß[ȣ)��9����!��3C��=j�s�$&�E99\2�q��Z�tk�n���lk{rŇ���n���c�W�ٺGb�n�������w�ğ
�H���E�u�{�c� ����=���a�C�M4 XۮW>L}q��M6�1��L�L�����t�U
��;�7uλ{�aT|�,���L6J/F�p#�{	X2��{Єi�$7����� �C�pL�����OCE��i}:у.�t���>9��F�b�Z)Gl��j�ﻟ(p���S�&��C���	��y ���h>�ࠃ9:%I
+ġan}��T���!�#���3��g����������wve�VVU��gc'�2
�$qw����0�׸.	4�|���kA�:0��f����[V�H1���"G�c��r�Onu�с�m�c�ی�^��1��nV쪦)2e�$5̒VZa�)��a6��`�+ N�:윥�9َ�9439�I��Bj�Ͳ��	&��X*�ɶP��������R�qn�l�H#�Uk�s��v���JhIG54���f�t�5��n�p�ɤî��Έ�n�8E�Ӆ8\�ۗ`G���)4�D#F}���������q�����HAJ �0�4���VM묊��خ��d�Gb��W�b�7}��q�$��3�a!�	�iА�;tte�|�!������n��CYٳ!e{ӻ�*��Yn�CF|�^�#ic���v�wp��\�6��l-��/�U�����i��Y��'C�l�Ä�/���cj	I8..ܺ%S�̅}�ćs�>(�	k^�����B|�1�<��`� �@hV ���vDxHЅWW1�Â���~ ��<I]@�c���ǁu�m8-5AM2g�"��J��g ���v-�s� ���xBnN�:��KƮ��sG�o�UVܒ����n,Gi�`B��u`Ϯ.�MV��D�Y6�Ӹ�7%�z1���bV�5p�������H0�uFp�A
���h�B��n�&�������ϫ��Gt�U�d��g��?d!:&|N��2z0���&E�=��Z��6����g��}�s�=���b"L�u��C)92��9#N���pk]��<6�$2���H6�V�Ɵl��W޻6a�!���c���&�(!T�L\8�����nIaI�.����y^(M�`?؏�fy�{�H2�Z6�����?&�1��6���C\={�fzz�v2�C���$��!�:A�V~��F�S�d��n���C�C41����=$��3
 �a@�\��c{)r�9�����4RGl���w!i��8\?;������JB�	���4=�8&�;�ك�E	���� d�h\\\�w]��c+ǳ�9�T�Tꝧ*5�5�{���L֣.G��4��}�3{��0���Ȋk�U����f{��΍�]�p�ND�7��;�������E?��ED_����y{rQ�E��ct�����>��њǻ�9�2���A:���t��E5�!���C)o�e=<?/�B�a���w���L�R��un��4|=6Op�o8$7�����ɧ�e�	���^Hg>���vЙ�������]�xk+�`�^���Z��0wOC�^�e�S�%0�@b�Z;�W�;�wн$����m��kG�7���7�Z�Ӆ��������ә�y�m]� WS��g��DF&�n8��ze�2��1��s��a!�G�^7���s��!3����Iƾ�R��Y���k�Cm�l`1���P�K����1
0�rq�w����uo#��к�F�%惣l�,�=�g�O��=b���Ue�7M��\K���!To���+�UI�^���c�`�Z"ő�5�4�L&�Q�7
{��~Z�$!��?Dόg4�2�1�;��e��>�6)�)n7i�Jv�^�A���ϥ�)*�yԻf�:$=��xG�_�d�� Ok7n�+�;2r"�a8��."X#�6��,W ÈN
n(�|4E+�x$=<�0t�bNBB��`P�d��e�lpj�K����o8�w8b.cr]��q���68S�udv��3�v��_r_<u��,�2��{����Y0p��7ηd]&�~��������f63�R\����k޺+~K}O�$�M�)�pv`��\�ڟzb>_���y	�,]g�����+�h���l�D���(P�>��{T5��C�ݕ���3�&�'C���v<��D����8D �7M�W,���|�a�$hA��0z3���P�U�B刡��#�߆�>!N$&c�-��i�m�TA�C"���E���F�qd�>K<#�h����������z;�Z>����=��'x�o�f��e��������S�cw�Ŋ�պ��O޽�h��"Rm<%$���?@�/g�N7�z�cۇ��P�,��Nwj���ݓ�jfFt5%�55��&Kl�����1˻0�=�G,q�SN�:ݔ���u�]`ҍ&�k7�M��qs�<��g�fOk��w��KJ:eu��9���"�DU��I\�IK�FSrJ�F�ؖ�5==sc�$�u�.�v�sy�S��N���K��}Zɓ���o�����.Ҩ�׀���5)���A" n��:16���1����3�t��ڧ��� ��}��fa���8�,�;�>�߉���/j��5�p�cLCi�������	S�i���N�;��:o�x��ve	��_�4�)� �Xc
!��xh�N����Dďa�k�tEX(y�L�'����*�)���GxW�aDCP�0�,�*�~�D����o�.'���H���x$2�W����F���!6ӈ �a ��ѵ&\d�`�P��_�*�M1~�c�öox��#;n7���j�!Bi�m& �Bξ���:�y#���k*�{o��n��GP�9Ƞ��,.iMz @��x��5��#y���+�WJ�v����C�n�h������Fcq��n�(�E!��|�Hg,���>��I�6����r�m��)�v������{-����OV̹�K����!���Y��y�ttES��k�)����j��LdG�� �H$���6g�q	����O�&�M�����;���9�N@H�U:�v��f�N�[T"���)�&]N�A����>�0'Ey���mD|�%7���@H3Y��@�k�_{�B٫�G���o>|o�Ɓ���m��az��JF�rD�
P�{�L����K�����k�s�$K��mU`��s�&��{dm��I!����߿�E�����E|B�bA���|4>Uc��}��tO�"M�I!�0C�$\cl�m��\sº%G.m�(�&�39lۭl�g��ˊ��d�wTQ,x�+��!���t��7��|ex�����f�:����;D���돡�)�Z&���'WG�@�c���"툞d'���������W&����PL1��o�� ��������l�?� yG�I��e��ǽ7�Wћ:�}�A�{��:f��]�9�"�s�Ӫ X�1V.�E�gO�I�R�V�SQ*�1��A�o�VVee�1��}�`0Ɵ��1�g{#2�1�m�c,t'�v�ن��`p�А��w� �N��a�WWb"w��h�a�C)� $F3�4H��Lv��f�, |����J�D������ �A ��~��>�zd�do�b��6s�*m���#�f���O%o#lEV�n��o3�~]�{�oZē3[v\3*~=��.�=8466&�8s��;��Hl�7mE�h�J(دu�l�� �HĔ?C��Ӧ}��r����D&�p{�*����C���eg>s�%�7�@� ���8<���/�}7U�6N��P�H��<~�А��u{ܹ)���2�	0a�({�=�8̎�u��01�xhZ2pc�w��c��[�x{�.7�ou<���/
��/uh[�˫?F��r"Dvu��De�[o�>�9�"6m��+E��q.b���������Ƹ���A0�&+^�w�"Eh��>�n����M����>O� ���/���?z��Ys�k�#��{$��ޞzA��5�ݳp;Ɗ��=��#�c��汮��WF[i!����Q��m�hm�z�ӿ�+�Y����3�8���/U�P�>�V�A�����L'���:ssuDs�In��Ē8o�6	�B�AS����?����J 4�I����P�0�D��'9����D#c���w�,��g� ��\ ���!A-��
����N��5��	C��hѲ�p��z���Fs�>�.a�MD<pJ4w��1u"s��8l	����i�k}:9�]=������S�����&�ظ�m�m�.�5��m��xq���	.�c�H� "iƀB5���ZkMh�ƫJV�5�jiU�m65clY5��RmmE�Q�[I�QmRm�6�b�6�Ѩ��mV6��cV�ɪ��TZբ��j��գl[m��kc[V��Q�Y-kVM��Rխ[�[%k4��[Xֲ��MV6�Smb�i6�6�6�-h�b����+E���m���5�m�h�Z����[[�V�Ze�Z�jekd�RjűV��%m�m�-�j�6���,�mcZ+b�l�ێ�kW&թ6�jڊ�5X�j+Z�j�j�m�mm�mUX�Vѭ��i��t��\���KmkEZ�ˊЩ�M�@]8� .��� ��Z�6�5Z�F֫�cZ�[[��km�m\5��ָkU��5Q���X�*�-�E�����*�[b�Qm�6�Ekq5X��)�ԥ����ڔ��wӗ��8�e]2t��*�ն�Y7]׼��]<v������WܮM~���\�C,�7י�w��Fu�󭭫m���|�ٮ�w_�m��m������l��U����]߻kqk��W��}��W�W��Ӗ�}�m�-�o���_?��r��.�W�m���ھ��q뫍/��{��)��Mu���Ys]��;�߽ۍ��[����Ʈ��黷J��[�SwU縶��k��_Fۿ5p���I	/ޭ5 $&$�\H�)4k�*L�Ih!���f� �&0h�%�h,c4a"ƈŘi$66,4��XH�f��2P�2b�b2i���bJ�QE��!)2`�10��2�X�`��i(1&*CQ!h�*(�&31I��%$&)�*1�Lز�!6*Mj4Q�HX�XI
�	�cE��Db�ш�fb�E`�5$��E�%��(1��f#�Ĕc�"�h��E��BJad,X��m$&,�E�س1)�"EF�%$)1�
d�c(��E&�4Ff�!��#%%& �b1l�(0bLh��l��jC!�H�A!�R%BbƌQD�Bh�Y(�FBA!EX��I���A�FB��c��#!���I�(4���Bf$T��cF(�%6)1�ĕfȘ�Q`����SLH�36bC ١I)	!�&)0����Ȥ�ƂD�dfQ#��b$Pə�L�Bc10�
bA����JYd&ja!)�`�����K1HHi,2d!�"Hi�(��Q�$�&2i�$�4Y(��2�$d�31��I�1$S3(�D�LĤd2	b�)��1I#4,��I��4I���ҊHLd�&)L���E&�)�$R(LL�D�4����H�IBF��i̘�$�1IB��"L&�ś"ME�$�3LRX�Ja
J20�,�&��4�ɡ�%#L�(ɊBɍ4$�����f4�dĆ��0�6LI�Sd$�I������&�fLѓ�(�Q&Ɠbe%���Ld�%���cIFLS(J*M���Œ2c%%(�b�$�d�R&i(��i�i
H�Œ�(T��4�&3#I�HdĖ&��b�H�S,Hi(�bSK	FHɌȐL&��(�"�L��M2)I���"X��ؓ�4��1�+A��lcj�h�ƪ�Qh�XԶګ+EX�kE��+b�5�TUX�5�UY5�b�Z�Ջ��6��E���U��ڋhڢ�[1�Z�+UDh�4TZ6����F�65���b+jKDkj�#E��b�kF�h�Qb�b�6�Z(����Eh�&ѴDmF��DmF��4D��X�1���5�TV�ch��,EF�Q�[�Ekk�2Qh�QQ�F�������clV�E�j6�}��ո�ڒ(֢ō��lERY)5��IX��6��(�#m���ѴZ5�j5�QY#h���6�6�cIj6�6�lF��Z4V55EE������,Qfk2�Q�hأ���(��jMbJ��-������̈�Z6KI(�%5EF�$���II���#cT�,TE�E�$�JKm&�kQ�Qi(�I$��TDmH�Y*(�RX�6�-$�,X�b"*H�Y*(��h��Dd��d�E�"1l���cb,RlE��$�d�Dh�mɴEEFJ�jH�,D�H��&�"��Ƣ-�DV1��Ԗ"�F��6Ƭh�QK65F�"���2أe���Ib5$��%�I(�d�"�Ql��DX�J#l�b�$b(��lM*f�",lh���I#DRj(�RE""�Dm%$��2�I�"I$�"�DcD���EX��e�I��,�ci(�*&E$�AY4DQDQX��آ�$I�JKF�DQL�E�$��S6"��F�F�&�5Q���4�%�I-�&T����F��KF�Ѵh�Z"-����Q%��F�#b(��lm$V1&JJ���#b6�&�Rh�d�DZ$�,m�,,�X��h��Qb�ɨ�X�kDDF�E����ň�b��M�IFƢ��F�5ERlQ�.��p�F�bH��cj(�"I+ID�h���Ѣ"�b��ƱQ��(�k����IQD���6�U�XɊ�ZԈ��IQ��m-��F�Mh�QlZ*���-I�Tb��%�*��ŋ2ɶ+E�j6��j"6�j6��h�VJ�X�D�kb�6,V(�5�ڋ�(ъ�+QDclZ5F�,���F�lZ*�m��6*$�Z$�,I�h��I�b+E�hڒ�KcZ5DY��5�#Tj"5lQ�lj66�m�[%lm��,QEX�$���Q�lF�EDX�F��F�V*6�(��6�؍�[&�Ƣ��m�[�i#X�Ŋ�h��mV�Xص���bKF1&�E���Ƭj+�ԛQY*�5F�m��j�lm���b4Z,mF�Q�J�h�hڋ��Z5Eb-��cTV6���E�,kƬ�Qb֊��X������$ر���%��V,���#X���j*��Q�bƨ�h�j"��bŌ��m$mU��E�[�����Tm���j6�h�6*M��I�lČ*���d���Ce0�M��l�(��	K�RL�d1�%0�K	�3Ja2�"���M�IA$�)	� ���	-�)�J	UD���X�����c���h�c$�XɌE�`�20c0�A%E&��4 ��#4�%�c$2mc"cS%4`�(�L��A`�QI��i���1�F2& ��0h�M�H��RTbɩ1EHc&1�c0��BAI3b�DfQE�T[���or��w��wƶ�����k���x�پ���۞�ޛ{\_g);m�������>���z�ڿ�寳�������xkkj�n7o�}Ws�ӵ��ލ��f�s��m���y���+~|�����w����_����C�W�����/����$���?D�Ё@
AV�^�|/?��n.�*��^��7�mm�m�+kj�o��<�ϫ��}��o�W+t�=[�~�$$	%�G�����҂�K���&�B@�LM_�MAB�8T6
4�� ����մ������Z�����qq.!���$	$�?(?a���]��k[V�sߓr�[�Rmj��m��u�o����x_&���E��u������]����n����}����m��ymڋy����onֶ���]��|+m�_��7v��y���۝��|7��|9ק*Y��^���^�����*	�~��v�b�E-��_�����pL���pxM~��0濐�HJ(�ê���x_��,e
#��8�Z�V6�Qm�ɛ�o���z�m�}-t����o���5�o<��k��ն�en
��[���	%�G��Ť�����X��_���-+-n�}۞�n����_���_m����������d�Mf���0�{~�Ae��������������                      ä���	��T��JRR�����D�@�� J�"�&�J��J
���3I������Ӯz�^���e�\f�����m���,vbu�� �v;zӲ;�Oz�ץ�ݮVtdm�68]��v�,u�ǣ(���@ ���*��H�{���<��WV��U�*\��ONʼ۶��u���j���]תO]ت�à�������tꪽ�Sr+�{�媝��՝�vչ�Wj�����R=r��k\��F��^  x��"RQ"�;��Λ����&�*�nYW[�S�^��]�ֻj�i�q�-Ps����.Z�M�x  c;�+�����|�s�W�榪��cmӺkm{k�Y{ԫ�=�];�N���n۶�ۛvԞzP��J�UR��oJr�"�v�Ю�uR�zS�y���U5q�te\��TW=�署���qj����
];{�Ӄ�ޏnw.�޲�yGvx���O^��z6�l{ K
P�I@c�^+��9<��oGH��;��t�3�]nî�#��K��ez��� 4���n����a�*k��7n�n�̦�Niݒ�0me}�
      0�IIT��hi�@�2@  fU@J*M� b@ @���R�jz��       '����	� i�	���2�F�d	��d�O �4hi�̉�A&����R0� � ��4�i�oG�.p赭jpu�(��Ei��ҩ�� ��DP- H"|���|lB�� @�"�e �cb�~'�#����3�}�3m<�Z�Ɇ�����L��X@�	,Q� @��r/@��(�n�EԀ��V�����U&$0��"�(�욡�ӧml���e���zJ��eT2��X�� �TQ�ݖxaX�ϡ�4q�8�,f���yS�O+ʅ�`�D$�������7����?�	��
�y��]�A�<I��/yd��f������}nʑ���z�wi�/;2;֣].n�[`ھ�0��xFn��ͮ[{S.jţ-7TSnv"��Wv�E�Ϻ�4�B�֭�Ƞ�,�NE���>y��M��{N!0\⒳$����כ7C=�'f�u<wd^�A��qM�Rtv��ď_,���}ܗ3ط��\�����D�C�p m��a�'F2��<%�v�jf5�i���m�>˸2���y����_e���ܻA���!�	����+�;�r�8���ރ�΋{Gxm��6����tYў&f�-� �oz��ܗ�]�$��R9��%���l[��y��6�fun	�f	��KDg,���Y��Z�8��8�S�:C��ؼ&�wv��������x]�x�ȷ���Ybͻ2�,��Y�uŪd���0�q=o����J,;��rv�J�����6�XH�O���ȝ��V��	+|pa�X���,��Ә��g�g5،Fu�/g`�p=�XF�ˌ<nw#t��w�ُ7o{{;&.\:�;��X�b�n�ᗺmm�y�0K��D��.c�u�.C��䰓�DR���>L[}�Հ���9�c�4�aɍ��a=.s:���x���&z�Y}9����K/lv�2�*��j�vK"wf�c�-H^��p�_Y;���i9�6�2���E��v�I5nv@[�$��9��l}�{��ˁK�^p/n՛�����}�t���4yӬ+�Y&�6ի� ���+�l{5��53ۓF �����V��k3�kl������s��;h�d_a�n	�����w<�E�4u�����Ŧ9�5`/Sm;����mv���=�޾�p��nG����w�9Ik�����j���dnB^�;�we�JM�巫�Z�}:u�נ�yvʙ����#�o�I����0j��V��[��0k�lp{Ü�u�o�݌��'��&.�͙��\�0,Ã�t-ZN��X1�ֺ�됥$�)M���>���Z�s�P���P8�x�i�7b4����,v��-6wJ����a�D��,�Yqm��Y|�{}�ApY'M�|ֻ�e�^���67�˼6�ɖR�T��F��S�Ρ�y��n;e)k���=���;�W����R- ��G(�`o_5����T���9��C6)-���{���$9�K,���z'!c�mF@V�/o�õ,,���MI����6�DK�=�Hh��G)�f�8��a�NnR��wp̝�&�]�9������}��m4�������՛[����ט�K37G1��F!���h�ݢ�=Y�/�"�X�}�掝�m�C�Vw|C��v�,�Z�H0�r���A�Q��i�x�`�ѵ����zѤ!/;���D!���ݡ.�@Oc+v�R�Z2��^c���",p68�R`w>db�pbOVn>�5k��{��Xq�滲Ӷ���g�	ܝ����8�xlǪ�օͽYm���wBT��-V��\�U����&iCs�K��xXwfr�/9�C�ãow��I�:8$����`N�E�ww��a垝x�����P����6�0I�Ļ�<�l���$3{]ȃ�;0�p�ܕ��_5q퉳1�XWGc�yi�0vD$��������sU��KK��φ2�dF\祌(�v�ݼ7� J�f�WcsVŴ��$	Ü�k��	�/!���#���h-���}�V[<xB1fv-,���;�K��1+����zc��r���8D՜�Z]���0�4�����S0.�h��O�1<��)b\o��!cb�ݩ�#\öӂ'��V��)j��[gU���Dš��d�2�kO6��qδ�7���-�0�|A�2��N��|t��,^g^�c���4f��1�׍��3����vzsvp[ow�Ɖ3:	�����9��z�!��V�؈x�w��i��ϱ������;x����Z˗�$��Z�h\���n\�ƴ�;���^�91���}hL۾���p�ם���bJfr�w.�3��,�R�#�Qs8V��2���2�q����Z:t޻ǅgf����Y"�%o]�z%������O�]�[ѝh���X�.܋v�'b��ٗ�ι�w�{�J�7mf�=vu��w�_Y.���y�r�[�Ne�x3/o u��ˬm�VI�d�W�7�Q��>7�sHԦ�k]�
)�ǝ��S�gja,�5�9V�p��ז��!����&Ej�	�ݶ��Ë]�Aɭv���xC�u	nR�н׺��II�4w:Y<��س7Ki�.�{�5vھ}�LȜ�y��a�祷Ǟ	��dњ���l��p�9�;w8-�����Iv�(�_bهz:���1�=2ٲmZ����h�ä���2[Ǣ�Y�ܱ#+x�i[��Y��Y�f-�|;;pE
��zzn;��oWkYyW�BdՉ͚������j\�1޶moYZ��-��"���͸MԽ=|"���5�Θs��K�wS;eݩQ[���0qjvs����M�M+Ә��;m�3�mn��'L��y������g��Z��s���1�{�`�����u�c35.:�dc_hX������M�f�����$//s�dS�G�N�IQ�n���I�t�"�U�A����z1C���D�۷�lü	�:�"Mɫ�=����0A�ڝ�j���,�+b	4y�����os�چv2v�w�m�P�}���#|�p��w�re�j�`q�֤�^�-<����H:�+[�#onm���D��|�d�&(�gfa*F�s]�*�V�{zLEǺ�"��܃;y����	��"\�����]��&e�s��l�I�\�ԑ��F�tb�Ј36!%���9ۘ��$��n�`�ы�$rO�a�PO.�gl7��-��g/wN�MpM���6tF�v޵{;�Q�N_��K��'�d�M�^d8����c�L��ce����h��;fA9]��2�3��1��a��/u��!�.-.b���Ih��B��q��S8&��_(���vIW2kP���v��1�8F�N�7��̬׸o ������;��R��𗉒/�N��F��!��妤'�����dP[O2��A�rqNg�^1���	���X�z�L:Υ��M�s/6�����G����juZ�r�620I�zu��N/�\'.Y�5]�s�2!;�]��W��m��k���{b����8�93qMج�fr�}�� ���"]�fB��7[��5�9ϖ�:��ˋ3:v�K��e�w_'�%�۝�)'s&��]�ܖ�9�:�����b+5GQ�����/\�{72n��2;��-nR{b�Z�B�Xw�"VZ���%�m;�`żT���nX�QvH���e���6Ⱥ��!=-�ok�1YxU�%%s�N�����;�},��-s��׹��j�����ď-VD�#��Z�v����7���^.�=�:A9�9�3l��ri��kz���3;v���xvf���	�l�L��bm�O{�c��5�z6���v��4�3,��h�֘v���dZ��-e�ovn���Moζu�/f�����m�aK��=�!��WZï7[A�EH��춝�^��Wۦi��d��۸�>���q�	1ͱ�.gLG��Ƿv���m���tv����D-!7�ݦсݺ�B���Ruv��fnf^X,)Q(�<��'t;�L�)���vw�>e䌭Nw�G"�ח
\ӎ�6�ձ�b$Z5�	�9��w���{��w0��ݚĹ{�rf��6��7{p�}���h�}M�[�k�����Y���rˍ�B�}��ļ�s��ؒ��z��69�3n�f�E�Fu�_b<0���ٗ7YG3�g�v:m��1	jSf��1A��r;˘8��<F��������#����?�
0!�C���l�̿Q�Cձ��SYCM�I8����[�pÞ��C"� �,� �8`��"1ٌ���j��¶��� K�]̴YLK˭�6�mt��#] �C��X͗T�[q2�X� �°�^5�v���q��K�Q�2ʮ�r���1�VӶl&.v�Z���h�DslkP-t�m2:�Ҷ��eVQjʚocm�>�[�D����>��,���#o&32�Ŧ����mh�դ���SfkH�)��ĪT0����R�J���x�L]Y��/���4[t�rk�4�D��z5�+*%��mu��S%֣�؆H
��č���p����.��0&�9��Ve*̸j�5Y��cpm7���K�>3��G�4� ���M41F����SG��B[�Ǝz�#BkK[m����g�kWι�!��G�43T 1�unfF�`F��í%�����)�'8Dl�SV��\jJ�3,���kYK(+Vj0�B��B�L2� �a�)�GS`��R��� �%�V355���,�q(YlW�aF�T0鱠�u��d�k��f�K.��j.l6��f�D��Y�sBj�KB�W�$��&Ԅ�ek���u��@-�`Yl.[m�]�d�[A�J�i7=���k�S���&[cYea�r:�jP�n�ċ�D�p8�;�[e!ai��ŬM����k��n5/[kbQ�ӱ�f����h�xj���T�t�]��Vf&�Rɘ
Z��t"���.�-ڰ��#rv͎[���Ź(�:���rX�c�8�$���e�#5�a�4���Q�ZƙՍ�+V�c[մI,ZZ��ځh1W �]F�8�H�M)K[*G�ͱ5��[����ҽ� �.lR��m�45de��ն*��t�2�t�.��fβ�I��j��e�X�ҪYz��nb`[�2�D�Ж��r�h$��Bet� �5���u��h��32�C��靚kY��W�c(��.1Gvte+����'+k�-5Xh�R9wJ�bcRf�-L��*������H]\��mU%���1��a�	�Ͷ]K��cBR��e����Ai]�j���ٰSxjhM6����gP�)N��40ˀ��)e�0K��׷a��P�X]�B4m[�����2�hYf��m�ݦQt2�`L�; �&�.�T1��cf�d��њ_R�f��CdR�+n���K�f��9��Є+t[�Tֱ�Vhlvo
+��pR��Y�.ጢ�AZ�(����[*µs�XCk�(��C�ժ7y,6��h\�mP��Vk
ۣn� ����CM���	l����aq)H��]lc�2�<�Ku�z�\�9�G�].&ٱ��m�JF"ֲ�O�x�jv�f��aDZ�ŷmŹ�@LP�h�*j�9a�a6�Lۆ%�m5�[��Q�F�p,JL���g`��0���\Z[���@���qK�
h�RЮ��14��f�V�,��B�S�BZʵ�,Kqz7fi�� �	������Kc
!,2�R��_KES�q��|����2k�+5Yu"c]�U*�)�f�1Xjl4P���MRɸ҄�4�b���Ѩ2�(:�0;�f�� YCY\���u�����X^ h`��X
�[4&�n���7�1��k���,qZ�\�d6���ʶ!�&;VقQin�3׆\K,v�.j�����BREe�i������W6�kP�uF�bm�H�m]�`Z&:�`͡���R�#�)i؃�ź�ҚX����,����A��lԊ��]�QdeMLѱ%Ƈb&y��{B�\�º]+-�����k,��P5Yi��4�[O'�M�ۨ�V%������b��xڬ3���)�KHv����ě6Q֐�T/j�܊Ao.f���Bx4�,�̵��Q��}Q�X����:\M*P̾4��]�̹ ���3�kLX��	Wo��&=nk����jk�J�"�Ki-
\��h��`[���3��mT.�\R����R;�Jfd�(lU�\�l�qRX��bly���hjG����|�Q�١E��9�rA�U���j���[E؂�^74��cZM
km��\Z+a�P�.�owX�^�eJ�mq���וG�7Vj��t`mv#�� A�����e�(4H7V��YMr7l��0X椢�.�jAf&h�.�R���s7Wu#�f8����˚Z4�C\ْ9��ĺ�RN�6̲�:ݣ`��[YS6a���ѧ^m2�+���*��Д�մ�Ү�m �BbmQ�W2�JMbDi(�Wh[R�M,f�0J�����6K�+��l��AuƖ�)Z5�3p�J� ԑ�m�ɔ�W����v��Mbe������.�S;lv�h�s���Y+��4HX�6�ZF�:Xq�J�MbkM���"���F��B��#�*�k��jJ��e9��d�&%3֣k�)�t�ne���{'j�&�D���!4�l�]�*3����D���`=��[.;e�	��f�׳4�����R
&r���ZB�3(g`6���f���W&�	EtFb�qqPu�	�l35&b�K�@�5Ԧ��%5�<[�Zs��VFP������XRVF6�	�Ȃh%���"�ٶ�ka@f(P�%oS2�v՗L�[��DbY,-������c�/�Z��n�UB��Z@�&a��EtH]K�	�����9-lPJ���^8_�[A�m��ME����Z�f�Iu
�n�+��U�	��9wRX�R-9�1�w����Δ��s4���R�a`����w����4
2cqZ�.��M�
��3��)5�W5e����q��5�;[L���2��m[��!�ڊe�mO�n�锤�&p��� j]]|k|��]�Ha`�]J�K3k��w.��5 �,.���H5�\�ZCj�к�Lݐ5��cڒ�v�KV���u��V���K^IV�7�� 
(Ѩe� ���͝ ���rp5Z�׮�5�ݧ���F�C�;v�(�A EI����pFš	bK)��OzO��w�O��ȼ6:��&&����r���[�3����Т��1��s�f ���`�Ҵ�SQP��E�Q�Y1�q Z3%���h��V����eH�c{ �YG]����B]���RS�
�`����l
i�mb�lkR>�l%˓kD#�-΍M�7Vݨr���M&�cY��;�a �x1J_��Z�X�F8.Q�nr1�����vU켦Ţ�P�"b���e��AbCYlslv�Aݰ\i0-eIRփ�&xJ�hW�uKe��*������p�B��!t��fC���i�kn	�]�#�h�G4󋉗c
�s�؍a�D3sq��Į�utS��iv{-�\����&�ڙ�
uu̳\�X���37dБ�,!D����\4�n�(�y��YYt�6��#,1!5���7!.��p�jϝL��]����<ɕ�-v��"An;Va����5���WT��l�|F�T����^J�2�q���%m�v�G���Š��Y�JH�����@eam�C��n���j�%%cR��B����maH&�m#5ѡ�l�E��F#}�����N��O;��o�3޲����6	A�۴�a�`�d��cP5a����]�v�s��b�Z��U6Xi�5&r:�q�Pa�#U�M��m,��h��e.H�U���@��WJ��G]�+�1���Ѱѕj-�YU��j�4�A&��(�O��cN��/��~�3�-L�g3��?��>�2�O�,����h H�$S7ۯV��o�C ���or�N�fb�^��\mI�{���ܼ̪�$Q$Pw����\R�<;����sُ0(p�*¨K_:��V �%��/�{��cr�U6���B�u��l�6��n�V����w��o����Go	�,�0��]ݐ�ۗ���M��mHdŻ��
�Q�h����Z�<�����On=����!���n�� ���9��9$q��#�Y�wN��� �E���fY�y�\��,F*	��4�����+�|�@0Ń֜�%#-.۴i�r1-A��_Z�Ӻwv�x]T��$,��V����n�9̞9I��C�k�7�^�MY,�D�RX��EQ���V����>��]�t�v��♓����D�c���ۻw�mʽS��O7�� R((��"(�	�1`������ghٞ`��		�Ć��y�6ٗ[pe�M8J-�E$�wݟ�u^yj�(�s�sO�F�·���{��s�~��F8�]�4b��#~;=��`�osK����F�C��:�';��}����&�14�$��XɌ�ٱ���ѓf`���rVo=�m�Vj�]�;�^ |�B(**"�H�$�"�=��U�m�i�o\���B �ܷ�Z��DR��ی�^q��5�BfT1��U��"Y�P>��,�7>�f��h����F0��7�[l�ۃ3�*�B�c�)���w��M�uu���λ�.z�-��7��8�(9��w|X��/�g��l���6�Q@����˪*4`����ۮ)Bƨ� ��Gq��f�O�-5���X�M�0�iP������b@���Z#5zmh4��P�2�v��`P��n�&*� v�f%e�d����XL�ڮ�%�fm6�D�%bÒhM�q`-Ұ�&�v��" ]F�v6ٌ���Y����$�AȂ���@ym���Ѻsx � ��n^^s�ֵz������/�z�p�s����BJ�$P!-v�81L|�E����߸wb;[ߗVՔ��	>TI�%w�;��k;F�T��&��>I8cMM���@]�L#Jb�,�$� Xs�sW�9ǜ�@�����j�|VXT�ڲ�MV\�&��h�A�Ԃ8"hF{>�<X<(t�������Y� ��h@A�)#h)�С0"���	����퓲��� iQ$N���w�ʐ��S!�w�Unn�׶��4�U �>�
2c)�^������@z-ni~���#�H�^z��H�)&M���b؋_:��Ut4m�`$
�v��2p�[�~^	�!��T�p���%I��ź���&�pD$���uˠ���P���e�h�2�n�UGBz�;�yg�큄!�UA�������LN8Y߸xU��{�ɘ��iD	P1�Jlh4����I6����������EF@X�_9��;�ۺ���a�w��o��:�F@Pb�P	�EW�w�h�nB��ԅ	��Gω0��"Iў������nݜ�  r���C��$�6T�Fk545�rb�h���۫nҮ�F�]��޳0�m  ��!;�{ڏFo���|��8�qH�����9Üਊ�E �������>� �'9xP}�û�F���Ac�\ÿ����Z' *����m�	���bu�z�E&�h���@��U�;��j)���#���߸w�d�!H�JB�%[��A����\.Ʌ�b��� �گvY���UU�쿐��j��t�~���EVz@&�Qb�u����}�v�UT}�,	8Q�=��fa��?
�&��a�����
F�C�w�w�����=���h�֒4��ف�SZ$���!!�&{�ں.�ղ�}�ss�P5h���VDB�'6(���
J���q�hj���i����\��&hk��GVlj�j�х�� ������t-���hA��L�3��#jh��+Y�d�&�ڥ�%�32�}�գ�|Qt�#Ce�ڔY��J��*X�@�Yt5R��f*1�s(�X �#A�t,U#�	P˺:x�$��
 � γ�g=�33�P
�f��e��e�ٟ<�UF,c'@�=�u�)�4X��/�(�e�x�z�y�R4(�4@�����r�#������ g�gw��O���A`��*H�����E��0C�;������P7kw����~����N�=��x��X�Δv��FmAb�FP���}_~��ӻ��SNOn?fϙnB�
�;Ah�Ѷ�W���}�W�dbY��R&#A �i$�)%�	b����ޞ]vB߹ͽ>�(�$o�7��*��[�j�s��n��'�<�ޖs4��	�2+��L2q\!��<x��lFƩ��y�DI�E�DJ�H�>s�g/�:F���o ({�w���\*���G�,�Ih�U@arSiǇe������F-��O^�67y~��w�����ciOUUA<�QC�����o�9���������vފ��{7� �&*w�% ���k��5�0����6Z6�{ɍgZ�s-+�G�K.)�ݬ��웚�ԝ��oV:�v �i���� �B���2���;u�;m')�gvӡ4���4���Ձ&��>(��[i|�I`�#m�Z���l��R��YΗ���]�vo)��ٚ�5&nzY���]j=Ku㞺ӱ�p��<��8��gsے��/h��T��r>ۣoG��n�+�:_!^�x��t)iI[ :����t�9;���W��{���uz������������z�k�)[�#'�`���6�Y,o�����3���� �b;��$���vT�1m
e�P��>���ȿ�������7���;7�d)������َ�p���D��O��,>Q�X��Q(��p����!j]�P��>�����EU00�&��1"��a�+Ϳ��]֮���sE5�e�,4��L6�mCB�mu�;=B�9}����f-��>(�TD�._E�����g
 j�6����RrG$�u�^ ~���e�)ª�o�{�(\6=�@�4(6��k�x�Ͼ�7sZ6��(ĩ�cu��??y�����%M,��BRi$��~?���+�C߿z�u���.�ᾴr?UP��1��$�J$:�v���ҩ�K��7lƜ���qE�.���xw�w\9����,a��a�$^﹯�j�NB�.��i�U
��/NOf3�$cIt=UKo�㽣v�� UÞ����r.z��p��Ԑ������$��}���{�}n��@>�\�5m�7��k�k|����; w�}����]]z��Q!��0�A�A�@��Q����+�4�jT�[��XT�0�s)Źq���95bbS����7iB�SZ��5��G�4%��*��_E� P֕BUu�m��m�0��"XQ��qilV�͚��elFݙ�@�`]���A%�b�y��Òx�`�r�BcE��%&��`J<g�����x=xӟ�n� i �j�o7�e����Ϝ�}w�k�Üy�d�i��s~~�aa�q�n)�:���Ƿng�=/�v-���|Ac<*�|�����XH {�<x�[��3�8Tk1JN8�hN_{�����@o�w`���q��+��,}T����Y��*���(db��,W[`U��Ô����4��@[�6��y�m` �P�i��FI��w�}�ʺ*�զ��|���vø����oK���H�-���;�V>��dy�� �AX *������]�:��'�J�{k���#d�٦��z����P�va��\))�p��U0;������s6�s��.J&�,F�&Kt\�X+��@S��[��6��}�z��d�0���p�%�p�q�� ����ۇ~�&�I���s��Ӯ��j]���3��<�ϵ�h"Q�"!���I�6�\v�뾾����V��M��ۻ�]]6eb��FHF�Yi6�����w}�P�v��n~8��MI P��$�@�}���t���k}�>9͟8R.A Z�)Ƴ14ήt�����&�j9gt�	�$�a�U'p���v^p��ǹ�c�G9��^U�C~�;��^}m�B�z�=�n?��f��[M�=�������C#U�N&��lk�=���Ÿ��%77��xw���?�{���U���%��p���V"��[���"q2 jH�F���[��he6��]��f���X���]YB��T�3o�o/:�ygh�Uݟw��
G&��v^xUJطf���kO�Q8�]�m����|�r�hƓn~s�S3L�,P$�cZ�����������>ޞvO��s�w����,3$&��ƛ��$C�{�p�o��7U��5�64B�	��d	"F32T�$4i&�1lL5�]��b�uf�28"�\�P����8�Ms)mŶT	��ą�q�c��D��i�8�[�Tm�V����qm��i�J��p�c-�r�z��bZS6X4�Y�l!&��51m�6�� ��n0�v�F�3�r��$*ZM���n�"Lc�\���?/Ke	 ���]�������;�D�WuN�{gd:[ �"�|���f��� �d����w���� I���{���m5���R��j�����Aw�ǻn�+1b3��&"N[�
���Gc7��$.tD��D
,Y	��[T
G�SZ�ZG]���B�D�f S�4ڎ ׏7�Y�7| ]��y���fwe�y��̾��X�b�X�L�J�c(�DED���������������9�Yt5r�5��z�{0�!b �1�d�ض4�m5�C��{ڏGw��q�Q�P�=���Y�«�wvK]��.S�ss���ù��;�@�h
�4H�j��q�%�[�g��	���n ݑkMX���ˉ�{6ի�m��7�7l|;�^�n��8F�:����{n�{�s�fsu�����j�o�='�lVM���8��Ŋ@I�?������~��;��HT^���v�U]h�6{�e�̸b2&�^xS]l�na�1����f��|��4��&\�Z�۫@%Z8)��M$l�̃��u��׻����tP"��y5����{:�>���sg�9H����I	PT��j�48j!�����{��v��K%0H�E���4bA�/�� 9n�y<:�P$qo�3�o{�>����\J#$1&�J6!,I�����I)@P�������9?�2�������=�p���TH&�A��X�|�}���vP؛e�.mY���f`�iWH��@����~��V��v#���gP��o}P�b���坣|*�wvC߽��LP�ch���}��D�r0e�UB(+��z��q�;�Ֆf��_q(��Q�(g�@�Hq{�g�G:���l�$n2���nfk��
�p�{����ŷ�)Z�����Y��ӊw�ۧ�.	r-���nu�zi�ݼ@с�I6)��_�̱��n�Wc\��f1.�k�4�z� �N��P��=KM�$M�=8�����'l��/��#��E��6od#c����Z�Nl�5D�"&d�v�KZ��ceq;����8O^��� �X>��R��[9[��,3��y���q���<�n4��(z�|�u�/vr�<��=�,`�^k0���F�I�ܞ��|�!�!�ƋJ�=V�������
�E�^͢�j�v�(���7�z���Y�t�{����"n[��-���[fґ�;N��x�~/�ڡ~<f�rY����c�[��V�X9�bcI���N�zM����;iz�C�zKx:����%�5�6�@�����+;����i�rm�ٗ0�ǋ�F��y!�^���GJg���sx5���4���:][Ss�灜���P��a��+�.qz���ܵ��uyg�f�Z(��KA8f�e�B$P���,�:����x�Oj�xv�������H]�{׫@�������[8��,��v����ݳK%��Z����7�����'�h뀔02P�v�ݥ��^e�
�U)/)���\i��a�`�0.�6(�ph��MA԰���nb��3J�\Bj��bM�D�m�0��W �m,�;)�qV�n�p�KİƆ%�@�����a�b]bKll`�P̵-�"\&nK+�ѷm����^f�4����KeeL�CYQ5�f�юuD�؛L"��B���Â	�M,e54Q�mt.��k),�.�L�+괙��)u3bG�u�
��mERSkR��ꀅ��5��blMH�wfiOfgYF�E��f$�Y�K.�`�3AR�h��l�K2�c��zu�3)
�L�GD�Mrm�6ٹ	ר<N%if�Ӊ����Mb]*$f�rM�uY�$��]FS;k4�+K�4��y4nК嵷D�y�����|�8��k��J띒)�ɖ�+�P%��f[���ڣ�����֚�Z��.ԆB¶���!4��h�S98�&5�D�H�;K�&�4��M�-�,�"- C75�XF`��62gx���n�Fk�r���1Ʃ
-Ⱥ��D���t����u��9k�YRĚ�Y�*7UTH�x�[Z��h�:���?��y�O3�Q�N��^3Q�T�-&%�[u�(�,aR�^r����R�C�.�����
Ԫ�tKl�tf�e�k	X3:ėkE�9n͇$��eIL�l�0HE��Xݭ��ۈB`�k`���%Vۛ�؛�]��-�i,��*�N�#��&h��]6�ʱ�g�7�e�g�%�D4��c�Xo+WՁ��nm����{�hϴl��Q4I�d�AQ��."	,"�#�����]���5����F�>�'r�p��o[I�c�<���ۛ�fK;U����芆FZ��Y��lX�@�w�i������8i~��bʀ�Ph���%��Fҍ!n(\q8��{5�s�c����{��3��q!�{��}��{��w�I��M
���(h� 	z�s��	&|7��g'���#�#��ja7J  ;��#���3��7ů�b)$[���MDР@��{!�ۗ������2#H�qZ�ƾF��V#ꮵ�f�E¤�M=��� }	 �$ H�At��6�[Y�N)ꭝ���s�;���HJAdFH�վ�7��$QE�"�"�ooڽQWW�u��:��1%��b��DH��M(b�I�	b�Lƿ�}�s��'�S�7��w����;;�� {����2�l	HJj�(z���}�>ѻ~Mm�,��#h�*:n�^ʰkSK)� �2�,����p��:��~��wv� 3�|e�j�j�9���w�� A��s�x'�|�z�oDP�
��a���u�Yi�����ϰg�u�\s�^v#&�_)�f�s\�C5N���*��1Ad��F4@���(�������u�2��U�^�Ek�����J%MF���_R����5�dY��
#K=�<hZ�^?���9��Վ��"\2�!�Z�-�3�|�o�<\�#;�R�^��!�z�0��:����ſ�ݷZ�>�ĭv�q�d����X�F�u��1�8q�DPO[~(��y�g����@�bA~"�P
�ީ�ɬ�l��+�=�pH����+��i����֬�t|u����CJ�t�ׄ3W��6�j��L �$�;�wkm?��V=L!�`Y�Othrץ"@����.e�֥q��h���k��È�V��m��r�"J���Wk`�6����*h!��.�R��E�����Z\���"l��f\�1(WZ��R��U1K���Y4[�i�3Y�rA`�����n �G���u�k���i�)����'�#z��_�Z�����w�1��k��\<G9��&ҍqʯܻ�8ӟ�Q�DQb�"6)-q_�sks� $P������YS΂9x��k·ݟ��m]�]nS��x�s�V8�J���5:��
�ރM����&�Q_�:D?U_}p�=Һ�f�*c��׳5��<D I�K����(�
_ő�>��0����T|hyy���W[�L�ښ}Q���Ԍ�|R7TVb�K�*�����*K��C\��0���+p~��4����ο��T�(�q��y�~�	R�3 H�%�BI)��!��N8�h��q���&��K��J�
��-�m�;P���bc5̣�=x�3�md$���+��K"�ݶ%W�4�߼�C�Ϗ"��}ᤨ"R]}@�wޮ%���J~m7���HE����L����4�OA��#.2�0���4��3++;Ko2�O;�bc�;B=d&�<���U����I���22���B�G3,���x�-���zY�:�����4/_�ۧWw�5�����(�P*�������y���Б!@4C��f��l�Cw�>��+n���������P|�?J
*����A�@�^�l�3u�~���}
*黺>�|�{�<��5��ÚdR$bOCD��V4�&^Pm�\���7�5O�P�������*���ҙEgz������E�$�QB�n&�K�rE���u��t��TB�w���ao l���q�{^�~O� �o���T�w��g�޾??�>��c@T���E�k�.�S��Y�~�s+M���v#�I��{�>�|�y���c�A��xx a���|�	�ԺG��t�s�i��N֊$Qb���x�}�y��fb�TU������e��|���f���k�%ko��B�����2����<E�l߇��Da��Q9$B�)�$�%^�� �*���>R�I��S��3�`��ɰPVATX�Zx�n�����z@�;��â�hk�3\�M?6��5;#3�J���5�4���f�Z���1/� ��=
��W]8�7��)��+ȕ����do�i}
pB�]���P �D�<w���Ot������߁7��ID��g��3J��6a��0	Y����W�&���\�j4�T���� i1��A��F��f%������ßV�U����E��1@����iºmq�s�W]�ʁa4b���f�`K��&��+�f�|��*)�ƕ�%Ȳ��Z����n]�f��j ��ԣ��έ#G3�#las�#��4Wh�K��٩7���!���31�Ў��{���>���0s+�����ʽ �X,��S#@��\WAd�р���O��g,���V�i]Y�d.��+��8�0������a���eEּL9��7_T)����x��C���pb��K��4�Q�]������"0A�2hb0b�����u��W?'���!o��KѤX�_�Y��μp����F�o>,�#�00��ܙi��?�%E!�q�+�a�k���;V�wnlM5hX��Ϗ�H�:���'L��d�i-��W3 �1������5�T����G��+�x>5��"�V��4�;�JꫪxB>�oQH������4��w��!w�A]���,�ͭz��]����P�PF���Q�^|x�c���zC?�ο�IsWw���6������
;}+�S�~`a�_��G�#���	�����!����.��0�v3��"��>"����g}��t�U۸as�^��J�[)�k"4uƓ^���s��7ke����q�L�w�i�Q�v�]z�>�͉ETcz���[�n{Ƶ�����Jq+<�0�@���U�=�b���%�j�/2�dG�Ÿ�M;#+Y�0�Z��r S�(A�,�N���,n��Y�iH"��]dea&ͣ>�����@� ��Sq9Q��Z/
A+8�����a�Ʊn�xK�j���ɧN��5-�p�AP+��wSSu��w�0��d��yz2�X�Ȥ��[2�����1Ch�O�)��gr�q@�f�6��0e���`ɕ�"�(�yi��"�˃�D�rI�,�R�Yp�H��ѹ��v�x�8%�l&�»���2�Ȏ����nFtܼD�ӏI��tԵv�1�-9f^颯C�����5�ݺ�J ���;p�M���܁cj��Z��;�+��������#M��00Ǡ}?�dҩ��U�Uv�W�����i�{�P��g���Z�N�6F=����%/Ƈ��@}��3dc�~�Z}ޔu������&�ﵯ;uZ�H4R��K4sX����yi�1A|to�^�V͇�W~�)%jCL�&�q�}����")4��A �^\#M���8�-�b��k�
��A���y\t�>o|h�S�3�m:�~��B�*8]՝6B�ޜ=�~,�:{��qӞ�G\,R"zkJAT�M_@/����Ԇ@U���,���w6���k�y��ZQ
��"!1�h�ͤP�c24M�T#4�@DF(2MZfy�a����N����/��u"p��L*��i�����w����~�),Z%Y*J�����=�u�Z��Uv��j�V�o"�F�h�Ό#3���N�u�w���V�SϤ����", �,����_�{��e&ݹ����&_��?I&l|l������,���PX��+ms+�%o*i�i���y�ɂ8����G���~#M�����gJ8���(����|�9~.H"���~�zG����μt��z��+M��w���Ac/�=�5t#��`ag�8� /y��� .{�E�̮%;Mא�`�1�foz���-�h��VYQ����S��X�BJ��l4����`�=a��f4�վU�� 1��]��K,Qi�	T�!T��X�@CV\ �59�h�6Q��ԕ��uı�*+�_�Q��|�V�����X�������2.Q"��U|�}V��-��K�t:N������^|�~u|��N��/�q�}���(�J�(��3�.�;���D�������������4e����ɏ}�i�Qרk��4��}�`(*0_�Lo�˅��c���:���)������������|x�6T�.��4ٛ�%爴�rǍ���qӴ���e���u:�V�S���u,�%�)A��Be��4�4����������>���R�1��.f��ٖ���1�y�I���/^��X(	�(=﫭&8�ݠ�N~�G���@?�����_�$�r�3��uq���Q)KE �(����qs�������Ǯ����><}GN�}ȧ�Kŕ�=gZC\�qҐ���#��w�j�>��|G#x��Z�9wVwB�Bw�u�w��L���n��D����|x�������j�<F��C���\Jx����m=�V3� �@!5�F�PT�H*ȌO��UP���e���6 ��qV���HP!7(��E�J��<l�@aeN�4�^_s⎑foA�߽��H�JA~"�u\$���_�Vx����C��F>��,��_��ڐȅ�?!�����ܝ`1H}߻�nk������h��F���5CeB^���9�8aN��l@�<M�����8���A��}����b'? y���5�F܊��~�N��Z�N�~M~�^0�eg��
��q��Ӂ���x�,����"���[=�����y�9��k5�3�H���K�j8ڀ���߾q������|x�7��B�xC8Fk����X`Qz����WXwXV8�~n��G�η�Cu�{�Z�����q-��S�ߐUcX��M�s�	��}��z��8l��t�>�k���ࡈ���Zc��z��9ޔu��Pj>�y�m��J����6�I|C?y	�#��xV0�aX�n�xA"	z S�Rw�?=�t�p��"K*3����߆Č�L�I�a12�]�e�q��k# chy��VW;z��1�S��WS%k*c�����#�2��{NZ�Zuq��Ս&ݹ�Pq��w��<�{��n��u�U������?2Dg��)Ĭ�M;l���|����f?{��+u�ݳ���6�X�D�+��|�ĳ;��g}��t�P��6��(^U�6�����ŭ��1Eb���V4�;s7^7:()!*u��x�o���4���(�H�aF$4~�����Uv�ʻ�H�\M*j�kD[knAI,E��,�C������ԔlX��ƈFB`�lZz�\[k\�c�)浰=��A���F�J,5ѫ),��T���mJd���QM0�[�fB]���F�m�[�%f�0�4�Y�i��d	�����O��g��ΐ�#��pz ������z|�q�dB��l��*�`�PV@�ϊ:D38�)���SZ�Z��>��@hH�I
�I��S�?&��x�9��Iz8��y�ŕ���I	i�6@^��}U�di��J�k��k�Դ����pYT�m�y����6��ab$QD` ������n�TU�;u�;g@�ץ"��e&��LRp'��Kb�6�Ё �:������%�����Z�Lv����!
��{��Yt��ۈ��%`q���ь��^�y�뽸[�������M(;o�RjI%�8a��~49p|x�6gFU�`�7߁n骶��q?Nò+_/�B���y1�V��;~|g�}`�3�,n���'7��q���, DD? DG(���q�dҕ�M�����~�_��m�����ù����
3q����m���#�`0˦�fe<���,>};_5���c��I���ϓ���m�g��rE
KY�x8��Y���g=�bcĭe7E"v�x�;sߢ�9q�Ƈ��ő��
#~Af��&I�K��h�"�QDQH��k�~�G�������m���t�7M���r��Pm�c��k�p�?wƇ.������tYeޯ���~����%��$R*g��r��QQ��U�]���N%���
y�+��]�o�Q.�nD{n.�r�m�Ŗ	�a]0���/�������������<x���co}Ҏ�C���۠�27?����}(3��gy����D]*�0�{O{�y����N�,_���~`~����tav�(�fi`@:������ăR��>!�����;���';��i���c
4�	�HEUX.W��ӛ��Ӫ�U�m�~y�&��="Q��^x�7�%���#���n�em)��7̩������)�D1hGD�I&@�U^�������f4�������So� �Da[��ۭ��mn�(��_w�5�D���Ͽ|��V��;~p�
2I�
�����=���n��|vʺ�j��1���~l��{���m���܆��s��ķ��a�G�+�x�?}��hr��	��4�}�~���"���2bA�^��@G����I�G����Q=_>O��څ9�+%k(�>:p��zx����	��?/�<\J�h�Ir�ɶ<������d;X���ґ4��p�/G���0�5Ý!�a�1��֐�\.kN�g�!�o��c�dیwP�,�����ݮ�3-����h%d+-HKB�y)���]�;K�n��U�1;�n�v{����w2��2���;� dx�v3v��ޱ8��s��^ �t:n��:��v�y���i�Җf��cv�T�]�o^o7�C�0gYM�N9�̭�mjs�Kgwb�5&�{��7wFR�v��zv��m�׊�m�ʰ /	�u�.o%�]FЩ- рA�/��k�eiBe��t��9+Z��ݬ�h���-�i}���LP&�%��	���Vʍ4Uک���8j�f��������d6�XiF�k�z���:�"�Wu��ڌ�h-�e!���ȎGi��z�AR�tСPY�����%�b̮Ҵ�R��Uq�6��6(����]j�\��Iaqf�5�TK�c��IL��E+zӘW8��ˊ8�A+fIM�=E�����G�Y�[ZKR�/,�����Ri�xm%��[
鶕T2nЈ(�а.�qI�e�Q�F�P3[�5���cYAVŎ��aX0�։-@3..3R@�m�Zҙ�]���y�g:̋3�0[��E���f�N�]�su(B�-����pt"�.u5Q�b%v_hV�6�.�|BV˽|.W+P��J�3�������Z�كL�d�H������]6��D�:l6Sa��Z��V�b�0��7BW0�Y�]�mKI�!ZL�(I�l�%س�u���e�����LX�0n�T�P��1�����0��dn��muV%4�6�� ۨMoaGX(�]7��������@(�[T2�X		rL���Ɩ�jVE�V�a�1d�Ջ��b�"�ƚ�3G�X{���~�|�xP�FP�@�6��t����4єA� ųA��.`�v�[�ĸ��F�m�<R��n����Y�!����%�ԛL��:�*�&tsV��b�`�	�Տ�`�Mf]X,Ճw^KX��ծ��\LY�q���%�p��0�Y�H%q���:�}y��/���QS���aG[}�<�{�ׯft�> ՟o�}�iHX��C>!�Α���`X,�E<��u�cf?00ß��C���>��~�⎑fgA�������	y׎�#}��crDYj_���~:t߼�������;���Z4ؤ�-�$�z�[Z�X�Hv�`ZMh*�E�i_{㍄�'t!�~xC8C�tO��dw��C�e��0��?���2V-�sB�i���#i-�����)C!��MX�}Aٟ��Yv�(�fi`p�{���#�}�1-���<~Mg��<���E �X�����I�%&���L�fR�4#A�O��V���P�Hk��|�u�}�s�(������7uf�گ�;z�o�논�+iN��"�<��E���p|h~���1��_���꫟@q�[�Y���9\t�"*ȱc|���1��UY�|���W�1q�0�y׎#���_���F3�������L�2&d��W.�Z�!��`��Yj��vNH�#+�!��|���}��[����:C�tN�G�w�!jIH_��{�L�Ħ �������m���0��^�3�a��n8��Ͽx>'^%k(��yRW���U#�Ph�Ad*�bk�z��~���n��ӛ���Uۯ��N�>��?�׽]z�6�^Y�y�ʰIP�\�\h��l�	bI!`���b�Aa��eq)�&�=�Z�j��^6��Һ�D;]+�S����6�W���z���߁O�2"���"����e�\�A����-2ؤJ_�"����3������μu�5�������Vݺ��m:KF1�ڤ""�((_^W�>m�x�������M��(C}������ؔ�v�Qv�x>�����{Һ�m��Y���12��Ɩ@]�J8E����L�Ё��`K��+��w�)5��ѫ����_VB�x~M(�&;�� �#N��08۟�Q׬fDW�W�>q6������de�&�0��X�86�$1f�lT[�a�Ѿ�{<�_6}��e��I��WX9�c��mC� 4	 �k��pF��<Y_��Y^�(�����=��<x���.�n
���ɬ��m"*�$S�a�u�'���{�� �~ }�߱�QF�����~��-��Z�����F����󫗋޽�;���#jIAQ��w��u��WkYktӪ>��sC�~`i�_�0��^�<D�����/���
$ �Q$))�$3h�b���$a/Y,���5�� 7ũ���˥k�m`g\��j5��j�
��v�si� ]�0��[,ɪ�1[չ�9�J��a# )���ݸ��cv�f�Z\�b��0�j�ьS;`ntlЌ�sHP�-��*�B��k3�⺈�K\-���J"�a�s���]���o>,�8gs�PMz�"(�4���=�NC"���kݬz�6�^\��9�ħ�Yʋ�Ӕ���wV���S��S����~c�W@Ჳ�Y�4�^�jw`m���U�1���&F�!�9XW����F	���e��T����?v��9��&���}��fe��߿1��{���O�7���g<!�#B�>&H�I!�R�]u��0\c��ՠ�$�6\�'O�D=���4<����|�����,��@@�W�vζ�����)���Q�,�x1zh�F� Pȉ��A&�F"QE"ɩ�����m:�Wj�����@"�5�?{ؑ�p2��Y:�z����h��=
��ϜM�]��߳�ޖ��֮��S� ��Ya�sqm�""�mz���M8�w�+�;�+M�:�W`�6�y��2��,x��=(�f�~��(,UH���]N��ک�ߓy��ǘ։,3k+�6FeD�.e�p�d1�`R�R�T>��ő���q�3�TN���Mh����W��Y�|�Q��wBo=?Q�H�Ή�i���a�±d�`�^�ǎ��?(�JB݁�eo�A�����H�y�B�������w�TYn�?2�����u
Q�Ȉ)\K�z�ü�cI�m�*t~{�y��~�0\�����,�OJ_�>�xC:C�tNF����_��|�_QqS�Q�^��H��s���Sfց��Ԍ_��f?00¯�0�� 5@�5_Pu~�fw���_�~�$�t}�ۏ�~��x���{|a��ƓoMw�`q�{���r@S<l��Ϗ���澾��ow�ħi\�E�n�AQ�&
3LAY4��Ow^�uM��U�~g�"H���"����EFH�C^*�&ߛ��ۧ�s�����K���3bd� )h�%414l	D��H8��|Q�,��|dN7A�_$�߿�~q+�S�ߓ^̾0��v��q�g����5��#6.-�ͱ�\$�ʐא�!*��I����O��w��q�"�z5?W���z�ow�Hg/���c����#�|Ƈ��c������
�Eۮ~�mx~��R@����Y���@����G\J�jc��׳/4%k��*�XM�;��5��Z���p�*2),q��A�;�J;�k�W�^|�m��\-�g�i���_u; �d�����m�{
��+z���e|�FBI�m"aL@JE
>���r��㞸��B���A���k��n��e0��f��6�����Kb�(W]	b�x�ڥ�[4.�n�%�,hgQB-���X�F�,&�T���t`��]�k�%�ͳy��r�ًl�sZe�^���(ʮ��
VX�6,UF�]��Hk��:|��$Xe���
{��bcĭeL}ki��i�-Ym��g�M�o�A�x�[{��>C^�u����7��M��U���v�)�Vr����R�$�i]��y�����2N�Y�,�Ƞ���Y^|�l��|� đ��+z0����t�3x��>#��Pt_���Ek�󍦿{��3�X�m߃_gh1���'�����-�{V9��ʹa�Wk��V�h�LыMT<}�q7@v��5~�{�S����6k�B:a�Q�������P8L��ӏ��Pm���QW���������Y���g���I�0� ��|Fתy��k=���"�$��jv�^��*��Lq�z����xCr9��d�?�^_#L~��g+�Nӗ�;&�U��*�~Mw���䀶��h|���z��F�+��Yv�(�fV})�l���1`�A�kq� M3jf��(�WkOơ� ��I�֑�S翼WSoR��1��k�����v��q���z�Uf���{��jI?#����ޯ6|F�҄;���KH��n����Ɠ��V0�aX��(�������Z�4�Tצ�#��Zޗ��f�W�v�@��+�����F$��!� q^%����[��Nv��k�����9�I���4,����x�%|�U� �'k�91��A5��mM�JqM�Зk�[e��ݯR�o,�k���%%�ϖw�l�N�1e��q�E�ݣ�Z[:��t5f%��7[��	J\ۺ��^a�e�D�C�:�K������!)�z��tگ�G��a�R�ڲ����b�K�i���C�ĉ���z�ݥԩ��;q��
H�a��5��̒۝w;�-�d��i��T�Y*G�!�! <�%��Xv�����ώ��y�x�Ĺ,�/�3'M�"A���x?���h�:s��a_�~� ,����$p��G��a�|]{���>n��3��}�Ɔ{г�
�~i8�����_=��<�{��n�2 c"�xH�X�Z^VO��Vb�(h��l�L&1�ʈL�!�"IH!BB���g�}<�,��ƾ �?��4ُ�a׫�2T���,ת�>�⎑foA����t�OI^:l���xL������ß��(H!jZ\ ��Z�la���Tb�뮟_�<�w�ׯo��>_2�
)Pg��3�l�D�do�P�D�4<����ez�z7#��%�6럻���̬t�>ox�)�p��Dz�� p^�rDL�&�P2��l�!m�6˫ݕ��AN#wP����M4;y�<�t�����J:��z�洵Wwz�H��B��8�녽�+�Nӗ�2GO#��~4?}�ˑG#�i�1����(�n������"���Uf,�e	2DT�^�t�3t���s�_�І����z��T���s/��C�P{�p�8�|��
�x3��hX��^�W_8�7]���o�ĭ��1�4�H���'a�3yQq�������3&���L� �,a�}��u�i5w�A���4��*LqFd�2Ǉ�L\��%�c+ب��ι�i�KÜ�X�T��)�!�B�=V��\fS:���d��(�sVl��5
�Q3�a���U�7�X�4��mE�m��.B��aR�V�3���2M��M@����|~#�����U��4��zQ�huR�c�����7A�~�<N�J�T�o��V~���y��D�2,�DTYtq���ʻ���k��5���ظ�\r��E����!���׉�̸z��V%<F��횲�/_E�I��WP�Vǈ�f=`a�_�0�����D�P���=O�<�+7?0���	�����W�M����Ɔ��(�`�
T]���F�B�yЮT�J��h�uu����}�Xco{�>CY���a���p$�=���PI	W����׼�7����`��Qf��IcV ��&�x�g�z��uҺ�v��9�*�Kh�F�h��5��
(�R8~9�Օ.�ob��_��v������P����z��E�^:l�~�?�FBw�C}�Ǚ �"�R+��y��cos�G^�����+��i��$B@Xj]}��p�_*vnUj�E��w��y��ұ��eq��P4�A)"�X��M'7s�h�tq0ڦ\x�Η��u��f6����N���Ƨ�'FC	F�������w��
���՝6B�ޜG�L�{]m8������h��@�$Q�2"�5��\����412'��?��!�פ<G�C�����x?���R)���7�N��w��U�`�u�G
8ox�)�����R�>�mĭv�]��\���&1i5]�����zx��s�Æo04��}�C̸�1�mz�m��\��tWJ�*�$q�p�c�d����>�B]/�>�C:GNtNG��9	Q���=^/�����Pm�_~�mu�/5|���hƱ����MhH(DT��c5����sv���W��S��V'^%k+�N�v��ݾ��r��0��r9q��:���ߋ��׻]z�6��/�C�KЈ1"�Sl%12	$�$����|C<F}�b	 Q�.��ɟ�U�������Ņ÷Һ����k*��7�J����+�Z"HrKT��@.��9@n�Fm�SE޾�oS��ҡO;�cS�`�'���ΰ�}Ӎ���l)~|Kю?{���t��P�{]}۞�z�q�����]��"����ߛ����&���*?�E'3
��+���(9tT���/>�Wm��_�[C����-�p��Ks�J�u��8a��R��E/�}T�J���B�w�֓�ܠ�n~�G^��.~���������F@�12͛!HH(d�UX1�/ν骲��u��F��!k�����f5�YU��s,Ҥ���B�!v�ԉ�W!krC��)K�_gn���ChW)��b�t �f��h�6j�ɤZ�B�h��J@�Ɨ�e�7�P�*`�v&!	fh�i6�ʮ.�@[ ���)A�Bw������3��߼�\#�bw��%$EI�<Y[��W~}�&R����2��M��`�f�hg�_:x���<3H��@�֭�J��_��:C���Ƣ�Gu�~_�}:ù�Ɠn��(8Ӳvw�>>|�kW�$FF��8x�1�҄?��8�t��t�F����i5��0���G�+ࢉr@��1��4����6��8��Y���g���H�"a�
%�bY�6[�f%PT��[�#h_���5���i��!{=4�����Æw?\l�|Q^q�>?�������Q&���s��㯻���Ȉ	"���(6}�zC<Fz�3����_&�F���C���8��e�u��Yǧ��NXw}��8��]NW�����S�ֱ<��z�N�~Mg�a���`O�WIQ�����H��������?��|
�4���{9��É�$*c4���d�ĤGکb�դB�)�N]#�@xQ��=���45x><F*kµB� s���Y��c���Ķ�҄�A�V+F4&FTĮ3Z ��+��^O8�꩎ߓ^̾3�#C���R5/���{��{�x���-e E)0EF�CA&d��?k�����?�;O�_{p�3�~�M�V��R�}#�n��4��k�3XV8�}� �t�Y���/�v���ﵯJ՚.��C++������5
s<�S���0᳔<�����2�M$E�L�`*�r2�tZ¬�vkً`�>��z��۶��m��+�>C^�y�a�g��!M�tz&��H*�#E����\�Ȭ���5c ��q/7SN�L�汆k
��#N��K��F�V��an��;8��p�S�aX��2��v^��U���v���_Xo�X�m�|��qMp�_�����͒�2Hh�d�DȄ�DY&���4�B������������p���#���i��z��3�TӶ���X�x��
ߨ�/�e6n�׎m.s5Ҥ�Z,(jEst���|������Ʌ_lg��|Q�,���3����8�����	<i]DI^�,��\�u�%h�j,[%F������Ɔw>0���7�`q���X^��n�O�_��{X�d���0�czPG����n�� �=���ƺտy����m����Mw��i�UAJ�_�g[C]��i��3�S�t�m���/~�?���8l���q�����at�g���j�E\�-�h��n���Q�+a�!��LCDଧl7=��t��e�K)LP����mAf	sR�cXr�s�:�����B���4ֺR�*bZ�c���:Od	-�s{2؅6�Ӯ3��Ӌ�kNl�B*��/n�]������-�����+9�;�r���zu{��;C��,/,�]�<u5��ݘG	n9�I{�w�.�.�K;��n�{#��Ω�y.絝z^��������7<��zg�jf[|�^f'Y����2[88�{���{�^vOg�h���ᲷҴl��j`2!����eKck���C��l��:bPzY�g��~�I�-��m�p[������B��iNƕp�eX�-�zU����+sb�16�#Z�
�v��3*XR��WM�%�]	�7`�X�5�[(��sS9�q��Ѡ[xH]F�ml����v�36˩�0aGd�f$�u�e��bP�)��ؔlh�f+�5��V��ZC4v�a�\(mf��{	�2ަԘ $�h�j+],Kq��M��U���ښ;�](�ö�k`��͂K����X&4#��03��0hV�Z͘Z���7gG�Ttqh������V�}�`�E��-��Z�,���GjML�u���(�Ml@�Mz�Q"�:�M�BQ�1���Jb���J�����d�H��W���q1o3U��-m0k*!nÄ�U�ɋ�*2�M�FZY��-l�R��Y�rG�z�Ά��b$vX˒k5�i�Fc8c��*��3e����^���pˬnV����\�ƶ�\2�z�m-[ ����JVWX���%�[�p!!nl��\�iI1G���y���1���T����R=�R9��t�]J�9�%}�Մ̩���1�%����mjGa�b���])��j|�}����SԵZ˥"�Օ�6\�Y��`cLi��5K����%`KL�%sv@�Zh�F����#m&ef�4R�z��RSK�a�b|)��E!�3�G�n3��<ͱfM�U p�9��=�p�.s�n`9l�ΰk3X�e˗dZ"�a����g�:�g����������
s|�%;M�dR ������,�]��&�������Ab�Ȥ`¡۲��8�����u��gC�s?0[��/�"���g��~#���:��[�|*�h��'m)Goޠ�ngZ�`0Qc~��i�z�����ǩ�W�p���f�Qz�����z���4��u�a�µ��t�6c��W��D.0����	�M�[Yr����kX�+Pt�_�6��+��T�6��T)��V\��i��[5���s{����@R

##�Ɠ���֛��h���Þ�c߁TQEcDX`T�����~�N�>��>C^�u������V�V[w���F,������w�TӶ����'�f�Һ�8�׏�{Vh������W����PЌ�`�s+8�7�*�>#������〹$��������7�X�j� �/�����(�������O6��WL]�Wh̫�
�kam�>�7���x�~����W��9�XH�Da�.�����b�*�c��A}��п���.C�_�ӆt`a�U���4�v�(�fit�����%F��|C_:����u��4F6�@�M�d�&��!��L$IAA�6hK��G���q�>���%�x��PX�t�#"����+�z��OzPgs^���ݒ����޿�lI5uT}�zW�ݼ����w_�Ͷ@�J8D3�a@�L��8 �P�3�^)\�j�սS����⺞q+]��ߓ\���O�k��6����
!
)"B �@�����zYp����G*���1���Q��������n��p���N =UJ� �����9t�G�x?�>?^CN�����6@ߢ�Ш�q'~=t(W�AU�F���g����:C\��U�]���_���0�r��IǍ�jx&�0V����|�����H§t��Q�����8��S5 ��d+BV8�.&It�eݎ��)�~��4��p�O�Eښh����߾~���be��(�EPP�y)�}�6���Y(�(��0����⎑�.�;���9���"	���u<�������Ԇ!#�4=�|Y�U-7�`q�߾||���ׯ���� �c���.��5.�=�zC8F�G��~�~4<����?��J	�8����,i�Y\t�-��S�ޗ�뉛,���QJa�Kd�e�Yg�/�ފ��(�X��nM6B��ڡ�j뙍�l	Fj1I�]pi�hBmFm�j �\:5�i����+cuM)p4�[f!ę�dn��ΆJ��-�aZ�i��6�Y��� �H�IJ2`l�����r2�l+[�5�w0pA4��f��6����Ϝ~Ms�o�r�"�5�E$$?H�}֓o��M1`1��,Ȍ�\n<�����=}�c��@7����u�\-����� 0R�;�Ɔ�?�aA fA~8F�3�� i����@�J8D=}��nڒ#_8�^�Sh�H?�~Ծq��_�,�C��x�����w��#N��04�cg�}E�wt|wd�J��W_8�n��y�W�t�y��wܯ��")4���}�4�c��fnW��+-քv��4b�ծ2\L$�����V;�dA����x�wA���6,��^�� ��>�+�I��7
{��bu�VUL���IX�5�x����da�6so�%�`}B����~y�������m�̹ٵ`�֤� ��y��x���"ԅtN�G~�|g����]z�~o.�m��ܳm�u�FA��" �~����5Km�ߝ>Koߚ�<�+> o�S��Y��4$�`(�(#$Y93�=��m�Z��e�\�#f[e�J�Uѫ���:(�^��f����*�AD�2���Mo�Pco}�=@^����3�(+����{�ʄ�%��q;ߪi�K=k;Һú�]z�~n�����ow�i�AI������[����߮q��%�$#2����b����)�6[����ꌃ{^>�J"���%z�|��9��#� ܾ47�� '���L��a�~h��5��R��ķݽ�j�����=�W��9�t���~�]a�aX�m�����E����ꪡX$�K-��\�6�J�굧E���jۭ�Hl�B)B%j���$��N����mw��N���Ǝ�n{�u:�s�����n�՝6B�ޛ�~ S  ;�ő����w~,q�P@t����h�S���¾��o�įI=Z$R7���M8�=����6�JC#���~`kn����!�r���R
($�/:�����,4I�) [�=�ιw����IM6/�a����Uj�}�Ɔ{�M�o2���9
d:�S�RII"�PQ��]{V�����u��g[M-�@�w�׌�޲ܮ[[j軧����Տ�&۬��#�ψgH�H�df�>X�	b�k�@1a!�U��|�~o�*�la Q��GH�;����M?B��ұ:�O�~!*��$D�	��s�?&���0�eci�}	5��u�V���Z�:��~h��w�ׯz��Goޔ!��3�d�>L�Ć]#�������J����|����r� ��PS[FZ!Ma�>;W;��,H4ٔ�u�����[lb�R�t"kA�эE�=�\V44������4���W,a�D��k^T��J�{%��6��\�]P#�t"R��l5�[��2RLRF�E����b��n��g^����\G̎��J9am`�e�jF+ɌL�V�j�>|�~Y��Ӡ�W���Z�N�~Mg����{��[w��p�$�m-�~�6�<�רk�P�>_#J���ϳ|4�� e��y{׼�k�ʹ�jH�fƛ��*�?&{�u�k
�o����$N?8?z��l��8��=(�fic¨ U~�~#�Hkθ�3�~0�	�]}�Ā�{��ӏ�h8ۙ�����B�J�(��H4�:��\�2_^mr�b�IY4m>����iM���R�\�h��e��Wz�Y���п=�=X~N�&f�i�I��X�5�c��X��� �J�>�m��Xa[��3X$��$C$�D��&�#h��)L4$�01�(�Ր$ץ�P��.�=��q�6<�N��]�W�眱P�@
������~�f�]���U
���~���l�����f2�"�l�r��sv����:���h��q� ��|��U�$H��ֳ��ʂ�t�+3]o�̴���xH�A8�A�
Bbk��6�A�Z�D��_'IM{����u���;���$�N9�=��mn��77VnCi 8� �(�D����q&�z����TO�P�l|���h|H�]�o28�-zm��D\4��Fkj�R�t��E���Nf鸛��|�|Y B��*O�����HI�������C��ua!�� �&��K<��s�=Kxa����i:�F���F;bŜ\�zvwDjc]�=��s�P*�rơ�KuMY����&�f��X��j���/p�j��՜�7v���.6h�ۄc{���˸��r�^�Y1d��n@�7���� �˫d%�Z�aSE�m�܏F��<ˎr��e����x��$YW�Q���!��V@Fo`�4�#I�c���e�<CЁ�X�Q��j%�DlB���2�Lj�pj�~�C��������>����{�F7,��À�P��d;�ݽ��*��������;� 4A� �FQ�9��z�EF�Xج�[�7�F�Z� �m�緘�_�[JD�r8�)��35k�p%���CJڢ��L�38@��;��ۏU  �����X��13���<(P{�;�ۇ=�|$�(x (���@ԍ7>}o��p��UP^����s��oT	9X�4a"=	�m�:�s�_/u�n�U����t�jj�UF��\m\زL5��㻎�yv�;�� -'�	'��%��Qa%�1*l�U�i4f�k6�J��=�W�W9���� Q�FMu�{���e���\Go�
��Y���<)�U 1�#�k�C��c�([&k9�[�KwNG�{F�p��_t~q�pǰ�����v�|(V����~k�rB�K׶_v�f��� �S2b\g\p�Q���&�fB0�)�O;��2�}��a&vb#��"� 0HŒ�ɚ)-��aPRAI $���g���`1ic��[+p��T<�-m���is���Wf&�j�X��V��vh|i�b[f�c-�R�iC���4���v����5u+�^���Э&S�����ת���nŕ`��vK���6�A6ͺ�;YU���	�n�{8��`�|t~v���UVC��#���q
8�d�݄��{����s���#(#"D-��EhwW{���`�*) �w��{p�巘� T&w���$�x�g\x�@���gs�1�/�7�כo7̶B��L�T��t���B ���sv��΄7������|��݆�"�k�%.6�Y��6;4���Ȃ��m������쒽��MU(E����^b�C'����箜;��?<��Q2�iL	 �e,E�>^y��iV@��j� ��k2����~P��aN;�O�:뙆szyϭ�c��T#��:z6�.y������{�̺�Z666��7ߝw�m�$�b ���z=IVV��������v��p���۵��#!)D����-mRX.8@�#ְ�m(�1�� Xսз�����x��V��m��������� $@P�`v1K�t�^w3o3u���M�U	�ڳ^Y� u|;����r^��N��x��s������L�N�����V�Fl��h�"h{���nT�{����P���_o��~'����s�j����W"�b1����Bp�F |����zoֶ����c�����f2#y�^�)Ѫ�s������O���G$JA������+h�(�kys��ز�3�B���R���e�,�������. Z�@��BiH(�@�1DY)E��0IL�D���
�R�If�`��F�㋁%�<9y~Z��"a�?q�s�f3����q
ꪦF�/�D�b�Q(�q4�.�J�$�3�R\��M�q�߸o�۟R��ݽ���Zߡ6���F�5D����}��Y{�/=�4o���n'��p�:=���x��[���P����_o����7�� r+����h�1X�5 [~����f��Y����x���mn��_�.��b!d�Q�Ê��n�
o1A���R��V�0�`Pŵf��eO�u�_fk�ل`��+��B�\̮Ź��Whv��)�	F.��5-\�B��\�ð�SK�A���],Q0KP���]	�\L;��Ya�7;�f1t�!t�V�B��P�3+\3A��}��Y�7N�ۏ����q!2fa�*�"����ـ�n�;�7ú�Q��s�{T���q�w��]�LL(!��sz�{��) �Uz�p唊I
`�W^��~kN[m��)�s�޷������SER
f�{��ow�C��#B��͠r��B�`�$��h*[��^�u]��{�;�F�&�J��q��~y�Ͼ�t"ؙ�X�1�2%Ϟw��;��v��ό���M���U�����Řm��~�����(�{�	�A&�sǞ}��|�j��D�	�h׳su]��~�9�D�c����/ue�
W��ZB��%�[4�b����6Zh!`�"1��)!�xg\x�췋=CL���A�"���QƲ�K���Ὀ��9����w�}mGrD�g{��^y矗�1���6#1L�RFi�IH��LiW���9��߼|��;�GV�ݛ��"��ŋP-5����k�%%U��n<v�췝�}qG�u��stn�wn�ћ�JSl������tm�۲E+��@.Eq7�1�c���{����HȻ�_us!��3���k;F�ѻv��"��D�F�K^�̆�"9��ṓ�㻈��7��ʐD$|hq ��E"(�!����_��n��3��ޏ	R&�j-��yB���Z�hѺ7n�_�x!1a��)�XF�-���P�� �S����{~�����S\�9��@�$)H	S!�v�n����{����N�p��ܲ��Ck;F�^i9�7�t���RTcY��3�|\�jd�V(�(RU�Ϯ��}N�����s7�B�D:j<�u�ν��wo7�k��Ι�f��	9�9zׄ��8Q^k�^�2���t���M�����u&
8�gI������N�$$�b�AE��!=���Y�D�"�{n�+r�e&�r˼����}2�7���#ק��=��G.sw�����:]t6���g�z	�Yz�2�V�k��/1�kK���مb/pc�9&3�3��7i��#7�Xl2���8���e���ňB/���S�ܼ��;	����gm�;4�ynj˾���&�V5=ܲp���x�M�X�w�˾�1��|un�o���5�2v���X�vOK�O�������N�����|Q=�(˳ ��a������i^H�[,���Ͻ��k���{�H�hu���xe���]�,�A��4���� p�R��掖�G_���{w �v��F�x��p�|6{A�b���o���%��\�p5�e燺��]�v��S���^7��v'#���^��׹��^�����y�l��޽^�w�����XFO��rWJ+m���*�q���l�9w��۽��H���-,>���ذN�Ǭ��g+��K��O�����6-+-CMUAl�ۅ��[V)2˴հ����,X�eڶ]d�����N�7.�k�e0��1+� ܚ+40�p�+����V2�Eс��0Z���le�Uf�혗���	P����E��cA��u�U˵YfQ�k[����%���6�Kc��٬�#`�f��tI��a���.�2�@�ܘ7[p�a�k�c�������]��t��v�'4����=v��f�롑�],3��Zfn�D���8.ݢ]2��4��y2(Kk�fӄPS6�᫮�*�2b]���W9c1t���əm�s602��3+3�������g�w��%�n�l݌�#Lh՗�t�Z1�w=�M�I��;9�fk�rL���v"��)j�4�:�l�c��Ѥ�%���P�rpJ����J�[iif��Z���Y�#`F6`�'�e�f��ڙ-t�u2�f�,Pm8]sr�9���TԬם���E.
��ciUꂑ�XƗ`�қ�!����\�0�)�m}X[0Xhek�u*�3P;`�[���B�E�Z]�r�	�-*�&�6���j�\��
���K�FQ��#��t�\P�SnK/����ǫ���]�J��L��;a&����s��V��0R&+(ֱ۫�t@�j;M���<강��ۦzܭ����VN[L�L�L&�Αf��xå0ķ3ku�M�ݜD���L�83����ƄR���؈Fmf�slĲĳ#H0�Tv���<߿�2��
�A *���fCh�����c�p޻x��[ �7/7��mD�[�؎�Þݽ�vhu5@�`��c[��Z��r|�DU`��EW�Ǽ{�춷^^b��N�fI0a�A�$>�����g���c��B&�
���1��ؖV�8i�k���b����c�qס���f��p�n���m�ԍNy���i2��ID�PDҙ�I�I�H(�4}��v��>�mf����D�A�[υ������	�Si�g9���\���UX0doW�S�#P�6�72`9������NM�I�t8�k�{��|{�wvY��&�E4t�M�V�@�����3Y�GUq�^�U޹�o|�F

D�&m��s�t�ݸrs)t"FL׋�p�a���ѻ��wp)#�!�v�}����lX��}��_q�،U
�KP�U\��{���z(�Q���/�e�+ǂ�g����(�EF:�=v�ܸs0�y�w>~{2)���wj�I��[���v1E��0�6��z�e�� �H��wd;ݷ������>$k��=v�AN�mn���x�Z��
��Zј���[@�U�H�,d�w� �Ȉ� Ϯ�v�{nb�["%�V���#�p�N�4j����0m4�FE�P<x	��j������q���Ǽ{����Yy�� �C&2oլ��\���-�ʸ��ٸ㨓���(�0��^{�ѻv^f3~�{�������g(��7ݸ{wG٩�b1|��=�3$�+BT�^8Ԗ, �L���V^�x2�D)�y𵝣t�ݺ�^Z3�u�ؕ�wpܹ�g�n��ߖ�ŀ�y��Z|�hZhi610̑�"�&�4�JD� ���X���X�T�_kWwUVR�Ez�Ҭ��aY�hɵ4(*f݈�B��
v�4&��F�!G����)��0��DQ��vcLG:�նb�K5��6�d,.%YF5�l6�dԍ��d�06�cK*S�3ZեE�Xj��	�S$��a.�t�F��D$o�k�y��~=ǻ�/8���҂�[���!��Ѻtn�>���WM7\Ӿ��RnVDd�"���}��5cMce�MQ$T��_h���σ��`.d;����w�(��	�Z���g/\&	/׶_r��W��Q B�5�o{���l2\�k�4mC���Vm��j�%�I���Fnc�Ż�#�+�_rP�!���+�����v�uݽ�}�֌a�Hu��kB ����&oo��lE�$Q�A�A �j��Ch疷�@�P����~��f����j7+M:�p�oO9���9��dX)�DsV����j�R8!,!�lV�wffR�V1Ś�扊k�xw�wvY٧/1�����[�;�F���ѝ����&��H$,U`��}����֮�w}xH$3Z"?_zk�ٜ�(�0X��)�#%2RE�'-̻y���8aww�U�_<�ݐT���{����;~�ɕ"FN[������H�b�W^�yk�2���Ӓ L"E��	ƌ�օ��#k@`��}ׯ6�+=�w0Y�@�(�S^<���-U^o3����n��3fp�c"Ȫm�|nbBMA��T� �@֗aȐ���x�Z��Ѻ7n�z�+�H����^�@m��r;�o9���\�GL���m��6�=�{�;���MB�d	P$�BC3hdrL���BU�5L|���N9y��� ��Ѿ��l�cc�,�}���ӽ���{:R��"�@dL�KIBH�X��Ti6X��\�fCC�Q�s�ow]���}����H:[��e�x�Z�oY2	"�#øg4h�4�Y��n3�~�u�H�T%���B0ȴD�*H� I�fL�%}��T�fk1u##6֨��B*��8��Ya+1LXkt2�C#�
�vn�vE��-�	�n0m���+e�(�Bë�$$n֕�Q�,q�f�ȴ�K�]%��3J	(L�-��a�F�&�6S0�sB�6���v�V�!rJ���Վ*�j;T&������;��E�۽�wy�2ą��s_{ü{�7�\�u�a��_��PTUQbł��y�u�[VsY�xs�9v^Z3���D�F�=�\aImK;pY�7qۇ;txn�d�/�e� , UDYy���9�ff�k����:�"͑�ffv�}�4��-�2$!���1�EN[���2��'Cۅ�ɨ��B9�V�X&����lR�HM�1�_z|��ˎ����S2���X�h���:lPU��,�E$3<��UzJ�{{U��Ǿ��{���N]f)�����mg�h��gӹ4ь������D$���9\���U��otn�s)��u���,�S!�-%�
��L��(�a��^� nn�ow��v�F̆(_�l�븉4AREk��z��)�IH�Y�Ԏ�k[�<�|�D��H���km����y�����u��8�a�y�n��gd�kn�ԙ��!1I�MKR;�eʌ��CJh*Y[i��`78�f��Xb�ѝ��I��A�Bu�K�wn�&�>�Af%<\���(�о�:te�N��Z"�u��*u�u[n�Lf�����/�t�k�r�䰷[zq��g/w[|�:���YXK���Ƿ0��i�Ҙ+/s:�ѝ�m��R����t^�� �u�t���4׍�t�_��;�z��.�Ν�V�N�^[ڄ�U�l.Z=����5|���!9!,�+XO%���ܢ������2�bT��v�b;nFt��z�?��?`����*3$c���p�n�n����8hD�d}�הA)hz��Y{�/1^d6��:�pB�$�ہWlf����˙Z��W$P���TM ���ў�x����a�RqH����"�UD�&,YD�扡U��H��}����v�ĵ�h���x�we��t���1fg[�#pHqn�����D!04�d����TFD
���_^��KT�"E�6Pq��[�+7F�#�p�n�ֺ$�3Dx�.%�Yŵ�vi��HNF\�9*r����p�;��e�5Ϸ�uU���w��e��F
�+	��*#Q����EE"�E�s��<9ϭ��o흹N&�Z"���g�l�r9��1E����dw�=�u��, $�$@�y�&���� ���R�Y���;�}[�� !X��FHd�de�i�����$L`,��9�aJ_Y���l�g%���"-�״�]�M-���XF�qc��+�8��V�5+6�0Iy���p�s.#TKc�V�Ԇv�lfG6h%�6+tI�k%�J��p�	�u�S`��7P8��5	K��	2���!8���cł,���s�^:շM��&,`�-��n<���m���4F�ui�{�3�t�8S����	UTMV����g3��w8Ғ$���^����a.�F��V�,�{_H��"a��v3{���G��� ��ɛ��hF�9�h2���"�զ r!#RF�l��w\=������y�����t��(�f�vB�X�R(������ozw���f��Af� u����ff/t�#WZ�s�w�9�`,U��QJ�$�Y{�{�1g8��9�w�t����R���}������"e���s��vr̖\$�#Q�[J}�s�n�9��� �H �	:L� �S6DE{�沭uM���Y�9���i��Bf�Ӿ;���}��۷����\d)�(�g3���Ih���L�E4���,d����)�cq�=������B9���2 ����hʹr33<q�˓Fn)b�L(�*��b�s�f;�����U�YE7IfƔ��#��n@˒���HL�Ĝ��R�Y��MQ$M���ǜ�)Fٶ-,f�w+�������gv3�#����v�T�,� ��C���dy�7F�oE����}�*��)y/Y
d�Q�KA���A$�	�x����HM�����5K07��燁O�!�d�f&�;�m�k��&n���F����F^�����ٽ᱂*���H���K]��!���I�M(f\Փ�y�
�F�N]��n��)y.�^��Y�BQg�������c9�;��FHr@�MP�EP�7��߳f�=Q#[�7�ݸ}�����^3�@�&�F3E�#2!ո��v�QõuWu�I�ɪ�aʤ��t�D���&�;bf�Z�Z��(\�l�t���1�)�5C�P�8+�f���u�V�Ƙm�: �*�-�ɠcZ6	Ir���҂�����j쮼���\M]ޮ��s�8���؈�+$@��Y*�*��AAHk���t��QD1wp�ѻh�f�82	� &�o�u���m�$/ǣ�,��wn݀��d���z��7l�������ݸ^��⤍0�׫tP ������G#���-DJ$�KQ������p�U�-�n� `�"�s�n�{���PdQ�?}������wþ{�|���CV^��������QV"��X��Jh�(��$���&1��(`�&��IhZ��Y��5n˟-��(��$w>�x�E��;F��EUF��i$UH:�.ڽk�ﹳ{�#�Y�7myj�$dȜ�(��/1K�g3���>I�9P�S��4a��f�srm��P�-����➖����}��}��j��!�DA&�۽���� rB�C����`3�1{}ژq��C���;`(��E���R�Di�n���U�|z4A5��9�-��E���e��ǋ�����j�J�t�`((3Xs7��O����mՒh`, ��E�/ǭo�M���&�f��"�!n�u)��L��=��I� � I$@q�܇}�y�iv�h9�wǆ�  ۲����}��"㉳>�9�7l,C� A� ��&]�ysa�k�G��tn�ݹ��
��~��$@�Y�,�qѻ�v^ʪ&�Ȉ((1�.���kE����4�u�MX�mVj�h��2�P��h����d�E�2,# ��$Q}��9�7m��IP@�Q��� ��g�n�ݹy����26��ڙ�� t�(����������";��x�E��Vn��ǯ̱�ZU�2�;���Z��呖]G#�T�uB2(�@ ���mR��?� @��G$pS��֦
P8BD PMp [��z�10t���-E dPT=�V�* 	r("Ƞ" �  6"�0� �Ȉ��b�� ��@PBPE/�3U��ն���\�)Hh� �����Y`���(�+�%j��$� ��`�pۏ��R�;����W� Ј�-T���DZ�x�Q��F�*�c��؂�7S(�F��UL��2���Q�RC���M��F�P>�]��l5�u3g�A��D>'B""�����R!� ���^��B���=�t�z��2�����Ե���:�)��}( �$u�O+X!?g�z���Sm���`���
��" ~�`���)�1��ԪL>�1���cC�)L���=�wf����!ME'�0��*QEI$!!#�aݿ4:`��� @��֬HR��z�iU^��D��5E2�l
gHQ/��"��vѹ=.w�P`Y?>N�{��Rrq�_������9��
^��Ǒ�~C���ݐI�	�gO#���!�>[2����D"}�ߺH}���C��gpp�!H �#�PLE9��[|���
]�9㰱��g�n�'ia���ל�sAO��_U���a�^A7�GqtC�S�������;�r�=�o� @�֏��І�B���G�Ҭ�dx�#�]Ӵ�kR�rS_�!�D�+���$� @�O���
E�ބF3��� r��>�1<�=������ԃa@�b�|ҕCa����Ӛ���q�!-D�1:pLE0����
%{zn�_D[�ȍ�x� ��R�SC�z��~�`�8 @�h@kp�d���O��d�@P=��(�;D��R�}e�fi�k�zM�̃�q`[
������q�;�0�������oM��@?����@ �o���� �S�S�ID<�D'�� @��.췩,�����c�y#7��x#y��/�3�r��<\�2������c�E.�$*%#������a�e6F�&��YIV,hrX�69��E.fq� E}Z�G!M�c�J�7jVl B+�0(��ρ�;�D7j�DS]#��(���X@��LUN�}�7���A" "������d�;�Ls��lL}�yd��y�>GA΃p�^�GI�,�*`n�jR�c��bͿ�|�EJT��D��{�6��]��rE8P��>�4